module heichips25_usb_cdc (clk,
    ena,
    rst_n,
    usb_dn_en_o,
    usb_dn_rx_i,
    usb_dn_tx_o,
    usb_dp_en_o,
    usb_dp_rx_i,
    usb_dp_tx_o,
    usb_dp_up_o,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 output usb_dn_en_o;
 input usb_dn_rx_i;
 output usb_dn_tx_o;
 output usb_dp_en_o;
 input usb_dp_rx_i;
 output usb_dp_tx_o;
 output usb_dp_up_o;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire net39;
 wire \u_usb_cdc.addr[0] ;
 wire \u_usb_cdc.addr[1] ;
 wire \u_usb_cdc.addr[2] ;
 wire \u_usb_cdc.addr[3] ;
 wire \u_usb_cdc.addr[4] ;
 wire \u_usb_cdc.addr[5] ;
 wire \u_usb_cdc.addr[6] ;
 wire \u_usb_cdc.bus_reset ;
 wire \u_usb_cdc.clk_cnt_q[0] ;
 wire \u_usb_cdc.clk_cnt_q[1] ;
 wire \u_usb_cdc.clk_gate_q ;
 wire \u_usb_cdc.configured_o ;
 wire \u_usb_cdc.ctrl_stall ;
 wire \u_usb_cdc.endp[0] ;
 wire \u_usb_cdc.endp[1] ;
 wire \u_usb_cdc.endp[2] ;
 wire \u_usb_cdc.endp[3] ;
 wire \u_usb_cdc.rstn ;
 wire \u_usb_cdc.rstn_sq[1] ;
 wire \u_usb_cdc.sie_in_data_ack ;
 wire \u_usb_cdc.sie_in_req ;
 wire \u_usb_cdc.sie_out_data[0] ;
 wire \u_usb_cdc.sie_out_data[1] ;
 wire \u_usb_cdc.sie_out_data[2] ;
 wire \u_usb_cdc.sie_out_data[3] ;
 wire \u_usb_cdc.sie_out_data[4] ;
 wire \u_usb_cdc.sie_out_data[5] ;
 wire \u_usb_cdc.sie_out_data[6] ;
 wire \u_usb_cdc.sie_out_data[7] ;
 wire \u_usb_cdc.sie_out_err ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[63] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[71] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[11] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[14] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[18] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[23] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[26] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[28] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[29] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[31] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[35] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[38] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[51] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[54] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[59] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[62] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[64] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[65] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[66] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[67] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[68] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[69] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[6] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[70] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[71] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[0] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[1] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[2] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[3] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[4] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[5] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[6] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.class_q ;
 wire \u_usb_cdc.u_ctrl_endp.dev_state_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ;
 wire \u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.in_dir_q ;
 wire \u_usb_cdc.u_ctrl_endp.in_endp_q ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[4] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.rec_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.rec_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[10] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[11] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[4] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[7] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[8] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[9] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[7] ;
 wire \u_usb_cdc.u_sie.addr_q[0] ;
 wire \u_usb_cdc.u_sie.addr_q[1] ;
 wire \u_usb_cdc.u_sie.addr_q[2] ;
 wire \u_usb_cdc.u_sie.addr_q[3] ;
 wire \u_usb_cdc.u_sie.addr_q[4] ;
 wire \u_usb_cdc.u_sie.addr_q[5] ;
 wire \u_usb_cdc.u_sie.addr_q[6] ;
 wire \u_usb_cdc.u_sie.crc16_q[0] ;
 wire \u_usb_cdc.u_sie.crc16_q[10] ;
 wire \u_usb_cdc.u_sie.crc16_q[11] ;
 wire \u_usb_cdc.u_sie.crc16_q[12] ;
 wire \u_usb_cdc.u_sie.crc16_q[13] ;
 wire \u_usb_cdc.u_sie.crc16_q[14] ;
 wire \u_usb_cdc.u_sie.crc16_q[15] ;
 wire \u_usb_cdc.u_sie.crc16_q[1] ;
 wire \u_usb_cdc.u_sie.crc16_q[2] ;
 wire \u_usb_cdc.u_sie.crc16_q[3] ;
 wire \u_usb_cdc.u_sie.crc16_q[4] ;
 wire \u_usb_cdc.u_sie.crc16_q[5] ;
 wire \u_usb_cdc.u_sie.crc16_q[6] ;
 wire \u_usb_cdc.u_sie.crc16_q[7] ;
 wire \u_usb_cdc.u_sie.crc16_q[8] ;
 wire \u_usb_cdc.u_sie.crc16_q[9] ;
 wire \u_usb_cdc.u_sie.data_q[0] ;
 wire \u_usb_cdc.u_sie.data_q[1] ;
 wire \u_usb_cdc.u_sie.data_q[2] ;
 wire \u_usb_cdc.u_sie.data_q[3] ;
 wire \u_usb_cdc.u_sie.data_q[4] ;
 wire \u_usb_cdc.u_sie.data_q[5] ;
 wire \u_usb_cdc.u_sie.data_q[6] ;
 wire \u_usb_cdc.u_sie.data_q[7] ;
 wire \u_usb_cdc.u_sie.delay_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.delay_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.delay_cnt_q[2] ;
 wire \u_usb_cdc.u_sie.in_byte_q[0] ;
 wire \u_usb_cdc.u_sie.in_byte_q[1] ;
 wire \u_usb_cdc.u_sie.in_byte_q[2] ;
 wire \u_usb_cdc.u_sie.in_byte_q[3] ;
 wire \u_usb_cdc.u_sie.in_toggle_q[0] ;
 wire \u_usb_cdc.u_sie.in_toggle_q[1] ;
 wire \u_usb_cdc.u_sie.in_toggle_q[2] ;
 wire \u_usb_cdc.u_sie.in_zlp_q[0] ;
 wire \u_usb_cdc.u_sie.in_zlp_q[1] ;
 wire \u_usb_cdc.u_sie.out_eop_q ;
 wire \u_usb_cdc.u_sie.out_toggle_q[0] ;
 wire \u_usb_cdc.u_sie.out_toggle_q[1] ;
 wire \u_usb_cdc.u_sie.phy_state_q[10] ;
 wire \u_usb_cdc.u_sie.phy_state_q[11] ;
 wire \u_usb_cdc.u_sie.phy_state_q[1] ;
 wire \u_usb_cdc.u_sie.phy_state_q[2] ;
 wire \u_usb_cdc.u_sie.phy_state_q[3] ;
 wire \u_usb_cdc.u_sie.phy_state_q[4] ;
 wire \u_usb_cdc.u_sie.phy_state_q[5] ;
 wire \u_usb_cdc.u_sie.phy_state_q[6] ;
 wire \u_usb_cdc.u_sie.phy_state_q[7] ;
 wire \u_usb_cdc.u_sie.phy_state_q[8] ;
 wire \u_usb_cdc.u_sie.phy_state_q[9] ;
 wire \u_usb_cdc.u_sie.pid_q[0] ;
 wire \u_usb_cdc.u_sie.pid_q[1] ;
 wire \u_usb_cdc.u_sie.pid_q[2] ;
 wire \u_usb_cdc.u_sie.pid_q[3] ;
 wire \u_usb_cdc.u_sie.rx_data[0] ;
 wire \u_usb_cdc.u_sie.rx_data[1] ;
 wire \u_usb_cdc.u_sie.rx_data[2] ;
 wire \u_usb_cdc.u_sie.rx_data[3] ;
 wire \u_usb_cdc.u_sie.rx_data[4] ;
 wire \u_usb_cdc.u_sie.rx_data[5] ;
 wire \u_usb_cdc.u_sie.rx_data[6] ;
 wire \u_usb_cdc.u_sie.rx_data[7] ;
 wire \u_usb_cdc.u_sie.rx_err ;
 wire \u_usb_cdc.u_sie.rx_valid ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_en_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_eop_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_err_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_valid_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.se0_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[5] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.state_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.state_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.state_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[5] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[6] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ;
 wire net33;
 wire net34;
 wire net35;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire clk_regs;
 wire net36;
 wire net37;
 wire net38;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net32;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_3_0__leaf_clk_regs;
 wire clknet_3_1__leaf_clk_regs;
 wire clknet_3_2__leaf_clk_regs;
 wire clknet_3_3__leaf_clk_regs;
 wire clknet_3_4__leaf_clk_regs;
 wire clknet_3_5__leaf_clk_regs;
 wire clknet_3_6__leaf_clk_regs;
 wire clknet_3_7__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire [0:0] \u_usb_cdc.bulk_out_nak ;
 wire [0:0] \u_usb_cdc.in_ready_o ;
 wire [0:0] \u_usb_cdc.out_valid_o ;

 sg13g2_inv_1 _2051_ (.VDD(VPWR),
    .Y(_1908_),
    .A(net481),
    .VSS(VGND));
 sg13g2_inv_1 _2052_ (.VDD(VPWR),
    .Y(_1909_),
    .A(net299),
    .VSS(VGND));
 sg13g2_inv_1 _2053_ (.VDD(VPWR),
    .Y(_1910_),
    .A(net764),
    .VSS(VGND));
 sg13g2_inv_1 _2054_ (.VDD(VPWR),
    .Y(_1911_),
    .A(net762),
    .VSS(VGND));
 sg13g2_inv_1 _2055_ (.VDD(VPWR),
    .Y(_1912_),
    .A(net760),
    .VSS(VGND));
 sg13g2_inv_4 _2056_ (.A(net761),
    .Y(_1913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2057_ (.A(net1019),
    .Y(_1914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2058_ (.A(net759),
    .Y(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2059_ (.VDD(VPWR),
    .Y(_1916_),
    .A(net757),
    .VSS(VGND));
 sg13g2_inv_4 _2060_ (.A(net758),
    .Y(_1917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2061_ (.VDD(VPWR),
    .Y(_1918_),
    .A(net1037),
    .VSS(VGND));
 sg13g2_inv_2 _2062_ (.Y(_1919_),
    .A(net843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2063_ (.VDD(VPWR),
    .Y(_1920_),
    .A(net836),
    .VSS(VGND));
 sg13g2_inv_1 _2064_ (.VDD(VPWR),
    .Y(_1921_),
    .A(net835),
    .VSS(VGND));
 sg13g2_inv_1 _2065_ (.VDD(VPWR),
    .Y(_1922_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ),
    .VSS(VGND));
 sg13g2_inv_4 _2066_ (.A(net797),
    .Y(_1923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2067_ (.Y(_1924_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2068_ (.Y(_1925_),
    .A(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2069_ (.VDD(VPWR),
    .Y(_1926_),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .VSS(VGND));
 sg13g2_inv_1 _2070_ (.VDD(VPWR),
    .Y(_1927_),
    .A(net959),
    .VSS(VGND));
 sg13g2_inv_1 _2071_ (.VDD(VPWR),
    .Y(_1928_),
    .A(net949),
    .VSS(VGND));
 sg13g2_inv_2 _2072_ (.Y(_1929_),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2073_ (.VDD(VPWR),
    .Y(_1930_),
    .A(net156),
    .VSS(VGND));
 sg13g2_inv_1 _2074_ (.VDD(VPWR),
    .Y(_1931_),
    .A(\u_usb_cdc.u_sie.out_eop_q ),
    .VSS(VGND));
 sg13g2_inv_1 _2075_ (.VDD(VPWR),
    .Y(_1932_),
    .A(\u_usb_cdc.u_sie.pid_q[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2076_ (.VDD(VPWR),
    .Y(_1933_),
    .A(\u_usb_cdc.u_sie.pid_q[1] ),
    .VSS(VGND));
 sg13g2_inv_2 _2077_ (.Y(_1934_),
    .A(net998),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2078_ (.VDD(VPWR),
    .Y(_1935_),
    .A(net1028),
    .VSS(VGND));
 sg13g2_inv_1 _2079_ (.VDD(VPWR),
    .Y(_1936_),
    .A(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2080_ (.VDD(VPWR),
    .Y(_1937_),
    .A(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2081_ (.VDD(VPWR),
    .Y(_1938_),
    .A(net794),
    .VSS(VGND));
 sg13g2_inv_4 _2082_ (.A(net744),
    .Y(_1939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2083_ (.Y(_1940_),
    .A(net851),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2084_ (.VDD(VPWR),
    .Y(_1941_),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2085_ (.VDD(VPWR),
    .Y(_1942_),
    .A(net1001),
    .VSS(VGND));
 sg13g2_inv_4 _2086_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .Y(_1943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2087_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .Y(_1944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2088_ (.VDD(VPWR),
    .Y(_1945_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2089_ (.VDD(VPWR),
    .Y(_1946_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _2090_ (.VDD(VPWR),
    .Y(_1947_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _2091_ (.VDD(VPWR),
    .Y(_1948_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2092_ (.VDD(VPWR),
    .Y(_1949_),
    .A(net209),
    .VSS(VGND));
 sg13g2_inv_1 _2093_ (.VDD(VPWR),
    .Y(_1950_),
    .A(net310),
    .VSS(VGND));
 sg13g2_inv_1 _2094_ (.VDD(VPWR),
    .Y(_1951_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ),
    .VSS(VGND));
 sg13g2_inv_2 _2095_ (.Y(_1952_),
    .A(net338),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2096_ (.VDD(VPWR),
    .Y(_1953_),
    .A(net928),
    .VSS(VGND));
 sg13g2_inv_1 _2097_ (.VDD(VPWR),
    .Y(_1954_),
    .A(net910),
    .VSS(VGND));
 sg13g2_inv_1 _2098_ (.VDD(VPWR),
    .Y(_1955_),
    .A(\u_usb_cdc.u_sie.crc16_q[13] ),
    .VSS(VGND));
 sg13g2_inv_1 _2099_ (.VDD(VPWR),
    .Y(_1956_),
    .A(net913),
    .VSS(VGND));
 sg13g2_inv_1 _2100_ (.VDD(VPWR),
    .Y(_1957_),
    .A(\u_usb_cdc.u_sie.crc16_q[11] ),
    .VSS(VGND));
 sg13g2_inv_1 _2101_ (.VDD(VPWR),
    .Y(_1958_),
    .A(\u_usb_cdc.u_sie.crc16_q[10] ),
    .VSS(VGND));
 sg13g2_inv_1 _2102_ (.VDD(VPWR),
    .Y(_1959_),
    .A(net888),
    .VSS(VGND));
 sg13g2_inv_1 _2103_ (.VDD(VPWR),
    .Y(_1960_),
    .A(\u_usb_cdc.u_sie.data_q[6] ),
    .VSS(VGND));
 sg13g2_inv_1 _2104_ (.VDD(VPWR),
    .Y(_1961_),
    .A(net915),
    .VSS(VGND));
 sg13g2_inv_2 _2105_ (.Y(_1962_),
    .A(net530),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2106_ (.VDD(VPWR),
    .Y(_1963_),
    .A(net932),
    .VSS(VGND));
 sg13g2_inv_1 _2107_ (.VDD(VPWR),
    .Y(_1964_),
    .A(net902),
    .VSS(VGND));
 sg13g2_inv_1 _2108_ (.VDD(VPWR),
    .Y(_1965_),
    .A(net854),
    .VSS(VGND));
 sg13g2_inv_2 _2109_ (.Y(_1966_),
    .A(net539),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2110_ (.VDD(VPWR),
    .Y(_1967_),
    .A(net973),
    .VSS(VGND));
 sg13g2_inv_2 _2111_ (.Y(_1968_),
    .A(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2112_ (.Y(_1969_),
    .A(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2113_ (.VDD(VPWR),
    .Y(_1970_),
    .A(net418),
    .VSS(VGND));
 sg13g2_inv_1 _2114_ (.VDD(VPWR),
    .Y(_1971_),
    .A(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .VSS(VGND));
 sg13g2_inv_2 _2115_ (.Y(_1972_),
    .A(net921),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2116_ (.VDD(VPWR),
    .Y(_1973_),
    .A(net301),
    .VSS(VGND));
 sg13g2_inv_2 _2117_ (.Y(_1974_),
    .A(net504),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2118_ (.VDD(VPWR),
    .Y(_1975_),
    .A(net961),
    .VSS(VGND));
 sg13g2_inv_1 _2119_ (.VDD(VPWR),
    .Y(_1976_),
    .A(net274),
    .VSS(VGND));
 sg13g2_inv_1 _2120_ (.VDD(VPWR),
    .Y(_1977_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ),
    .VSS(VGND));
 sg13g2_inv_2 _2121_ (.Y(_1978_),
    .A(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2122_ (.VDD(VPWR),
    .Y(_1979_),
    .A(net924),
    .VSS(VGND));
 sg13g2_inv_1 _2123_ (.VDD(VPWR),
    .Y(_1980_),
    .A(net828),
    .VSS(VGND));
 sg13g2_inv_1 _2124_ (.VDD(VPWR),
    .Y(_1981_),
    .A(net826),
    .VSS(VGND));
 sg13g2_inv_1 _2125_ (.VDD(VPWR),
    .Y(_1982_),
    .A(net812),
    .VSS(VGND));
 sg13g2_inv_4 _2126_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .Y(_1983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2127_ (.VDD(VPWR),
    .Y(_1984_),
    .A(net1003),
    .VSS(VGND));
 sg13g2_inv_1 _2128_ (.VDD(VPWR),
    .Y(_1985_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _2129_ (.VDD(VPWR),
    .Y(_1986_),
    .A(net575),
    .VSS(VGND));
 sg13g2_inv_1 _2130_ (.VDD(VPWR),
    .Y(_0039_),
    .A(net49),
    .VSS(VGND));
 sg13g2_inv_1 _2131_ (.VDD(VPWR),
    .Y(_1987_),
    .A(net486),
    .VSS(VGND));
 sg13g2_inv_1 _2132_ (.VDD(VPWR),
    .Y(_1988_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ),
    .VSS(VGND));
 sg13g2_inv_1 _2133_ (.VDD(VPWR),
    .Y(_1989_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ),
    .VSS(VGND));
 sg13g2_inv_1 _2134_ (.VDD(VPWR),
    .Y(_1990_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ),
    .VSS(VGND));
 sg13g2_inv_1 _2135_ (.VDD(VPWR),
    .Y(_1991_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .VSS(VGND));
 sg13g2_inv_1 _2136_ (.VDD(VPWR),
    .Y(_1992_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ),
    .VSS(VGND));
 sg13g2_inv_1 _2137_ (.VDD(VPWR),
    .Y(_1993_),
    .A(net991),
    .VSS(VGND));
 sg13g2_inv_1 _2138_ (.VDD(VPWR),
    .Y(_1994_),
    .A(net383),
    .VSS(VGND));
 sg13g2_inv_1 _2139_ (.VDD(VPWR),
    .Y(_1995_),
    .A(net290),
    .VSS(VGND));
 sg13g2_inv_1 _2140_ (.VDD(VPWR),
    .Y(_1996_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[11] ),
    .VSS(VGND));
 sg13g2_inv_1 _2141_ (.VDD(VPWR),
    .Y(_1997_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ),
    .VSS(VGND));
 sg13g2_inv_1 _2142_ (.VDD(VPWR),
    .Y(_1998_),
    .A(net280),
    .VSS(VGND));
 sg13g2_inv_1 _2143_ (.VDD(VPWR),
    .Y(_1999_),
    .A(net272),
    .VSS(VGND));
 sg13g2_inv_1 _2144_ (.VDD(VPWR),
    .Y(_2000_),
    .A(net222),
    .VSS(VGND));
 sg13g2_inv_1 _2145_ (.VDD(VPWR),
    .Y(_2001_),
    .A(net372),
    .VSS(VGND));
 sg13g2_inv_1 _2146_ (.VDD(VPWR),
    .Y(_2002_),
    .A(net370),
    .VSS(VGND));
 sg13g2_inv_1 _2147_ (.VDD(VPWR),
    .Y(_2003_),
    .A(net374),
    .VSS(VGND));
 sg13g2_inv_1 _2148_ (.VDD(VPWR),
    .Y(_2004_),
    .A(net387),
    .VSS(VGND));
 sg13g2_inv_1 _2149_ (.VDD(VPWR),
    .Y(_2005_),
    .A(net938),
    .VSS(VGND));
 sg13g2_inv_1 _2150_ (.VDD(VPWR),
    .Y(_2006_),
    .A(net174),
    .VSS(VGND));
 sg13g2_inv_1 _2151_ (.VDD(VPWR),
    .Y(_2007_),
    .A(net368),
    .VSS(VGND));
 sg13g2_inv_1 _2152_ (.VDD(VPWR),
    .Y(_2008_),
    .A(net296),
    .VSS(VGND));
 sg13g2_inv_1 _2153_ (.VDD(VPWR),
    .Y(_2009_),
    .A(net259),
    .VSS(VGND));
 sg13g2_inv_1 _2154_ (.VDD(VPWR),
    .Y(_2010_),
    .A(net23),
    .VSS(VGND));
 sg13g2_inv_1 _2155_ (.VDD(VPWR),
    .Y(_2011_),
    .A(net244),
    .VSS(VGND));
 sg13g2_inv_1 _2156_ (.VDD(VPWR),
    .Y(_2012_),
    .A(net294),
    .VSS(VGND));
 sg13g2_inv_1 _2157_ (.VDD(VPWR),
    .Y(_2013_),
    .A(net264),
    .VSS(VGND));
 sg13g2_or2_1 _2158_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2014_),
    .B(\u_usb_cdc.endp[2] ),
    .A(\u_usb_cdc.endp[3] ));
 sg13g2_nor3_2 _2159_ (.A(net995),
    .B(net971),
    .C(net972),
    .Y(_2015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2160_ (.A(net768),
    .B(\u_usb_cdc.endp[3] ),
    .C(\u_usb_cdc.endp[2] ),
    .Y(_2016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2161_ (.A(net710),
    .B(_2016_),
    .Y(_2017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2162_ (.B1(net847),
    .VDD(VPWR),
    .Y(_2018_),
    .VSS(VGND),
    .A1(net710),
    .A2(_2016_));
 sg13g2_nor4_1 _2163_ (.A(net845),
    .B(net842),
    .C(net836),
    .D(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .Y(_2019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2164_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net754),
    .Y(_2020_),
    .A2(_2019_),
    .A1(_2018_));
 sg13g2_nand3b_1 _2165_ (.B(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .C(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ),
    .Y(_2021_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ));
 sg13g2_inv_2 _2166_ (.Y(_2022_),
    .A(_2021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2167_ (.A(net717),
    .B(_2022_),
    .Y(_2023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2168_ (.Y(_2024_),
    .A(net747),
    .B(_2021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2169_ (.Y(_2025_),
    .A(net626),
    .B(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _2170_ (.X(_2026_),
    .A(net1009),
    .B(_0059_),
    .C(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2171_ (.B(_0059_),
    .C(_0058_),
    .A(_0060_),
    .Y(_2027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2172_ (.A(net626),
    .B(_2027_),
    .Y(_2028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2173_ (.Y(_2029_),
    .B1(_2028_),
    .B2(net872),
    .A2(net709),
    .A1(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2174_ (.A(net643),
    .B(net873),
    .Y(_2030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2175_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2007_),
    .A2(_2025_),
    .Y(_0066_),
    .B1(_2030_));
 sg13g2_nand2_1 _2176_ (.Y(_0065_),
    .A(net717),
    .B(_2006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2177_ (.Y(_2031_),
    .A(_1943_),
    .B(net553),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2178_ (.B1(_2031_),
    .VDD(VPWR),
    .Y(_2032_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .A2(_1945_));
 sg13g2_nor2_1 _2179_ (.A(_1944_),
    .B(net556),
    .Y(_2033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2180_ (.A(_2032_),
    .B(_2033_),
    .Y(_2034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2181_ (.B1(_2034_),
    .VDD(VPWR),
    .Y(_2035_),
    .VSS(VGND),
    .A1(_1943_),
    .A2(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ));
 sg13g2_nor2_2 _2182_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .Y(_2036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2183_ (.Y(_2037_),
    .A(_1943_),
    .B(_1944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2184_ (.Y(_2038_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2185_ (.B(_2037_),
    .C(_2038_),
    .A(_2035_),
    .Y(_2039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2186_ (.A(net567),
    .B_N(net53),
    .Y(_2040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2187_ (.Y(_2041_),
    .B(net53),
    .A_N(net567),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2188_ (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .B(_2040_),
    .X(_2042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2189_ (.Y(_2043_),
    .A(net976),
    .B(_2040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2190_ (.Y(_2044_),
    .A(net961),
    .B(_2042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2191_ (.A(_1944_),
    .B(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .C(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ),
    .D(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ),
    .Y(_2045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2192_ (.A(net310),
    .B(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ),
    .Y(_2046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2193_ (.B(_1943_),
    .C(_2045_),
    .A(_0056_),
    .Y(_2047_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2046_));
 sg13g2_nand4_1 _2194_ (.B(_2039_),
    .C(_2042_),
    .A(net961),
    .Y(_2048_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2047_));
 sg13g2_nand4_1 _2195_ (.B(_1944_),
    .C(net314),
    .A(net1022),
    .Y(_2049_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2042_));
 sg13g2_nand2b_1 _2196_ (.Y(_0429_),
    .B(_2033_),
    .A_N(_2031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2197_ (.Y(_0430_),
    .B(_0429_),
    .A_N(net990),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2198_ (.Y(_0431_),
    .A(net990),
    .B(net707),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2199_ (.B1(_0431_),
    .VDD(VPWR),
    .Y(_0432_),
    .VSS(VGND),
    .A1(net572),
    .A2(_2043_));
 sg13g2_and4_1 _2200_ (.A(_2048_),
    .B(_2049_),
    .C(_0430_),
    .D(_0432_),
    .X(_0064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2201_ (.Y(_0433_),
    .A(net626),
    .B(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2202_ (.Y(_0434_),
    .A(_1921_),
    .B(net368),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2203_ (.A(_2022_),
    .B(_0433_),
    .C(_0434_),
    .Y(_0435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2204_ (.A(net751),
    .B(net753),
    .C(net465),
    .Y(_0436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2205_ (.VDD(VPWR),
    .Y(_0437_),
    .A(_0436_),
    .VSS(VGND));
 sg13g2_nand2b_1 _2206_ (.Y(_0438_),
    .B(_0436_),
    .A_N(_0435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2207_ (.A(net745),
    .B(_0438_),
    .X(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2208_ (.Y(_0440_),
    .A(net745),
    .B(_0438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2209_ (.Y(_0441_),
    .B(net838),
    .A_N(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2210_ (.Y(_0442_),
    .A(net759),
    .B(\u_usb_cdc.addr[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2211_ (.Y(_0443_),
    .A(net758),
    .B(\u_usb_cdc.addr[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2212_ (.B(\u_usb_cdc.addr[3] ),
    .A(net760),
    .X(_0444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2213_ (.Y(_0445_),
    .A(net763),
    .B(\u_usb_cdc.addr[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2214_ (.B(\u_usb_cdc.addr[1] ),
    .A(net762),
    .X(_0446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2215_ (.B(\u_usb_cdc.addr[2] ),
    .A(net761),
    .X(_0447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2216_ (.B(\u_usb_cdc.addr[5] ),
    .A(\u_usb_cdc.sie_out_data[5] ),
    .X(_0448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2217_ (.A(_0444_),
    .B(_0446_),
    .C(_0447_),
    .D(_0448_),
    .Y(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2218_ (.B(_0443_),
    .C(_0445_),
    .A(_0442_),
    .Y(_0450_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0449_));
 sg13g2_nor2_2 _2219_ (.A(_1932_),
    .B(net944),
    .Y(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2220_ (.Y(_0452_),
    .A(\u_usb_cdc.u_sie.pid_q[3] ),
    .B(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2221_ (.A(net998),
    .B(_0450_),
    .C(_0452_),
    .X(_0453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2222_ (.A(_1934_),
    .B(net1028),
    .Y(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2223_ (.Y(_0455_),
    .A(_0451_),
    .B(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2224_ (.B(\u_usb_cdc.sie_out_data[5] ),
    .A(net761),
    .X(_0456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2225_ (.B(net767),
    .A(net760),
    .X(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2226_ (.Y(_0458_),
    .A(_0456_),
    .B(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2227_ (.Y(_0459_),
    .A(net763),
    .B(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2228_ (.Y(_0460_),
    .A(net760),
    .B(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2229_ (.Y(_0461_),
    .A(_0459_),
    .B(_0460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2230_ (.B(_0461_),
    .A(_0458_),
    .X(_0462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2231_ (.Y(_0463_),
    .A(\u_usb_cdc.u_sie.data_q[3] ),
    .B(_0462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2232_ (.B(net759),
    .A(net762),
    .X(_0464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2233_ (.B(_0464_),
    .A(net766),
    .X(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2234_ (.Y(_0466_),
    .A(_0461_),
    .B(_0465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2235_ (.Y(_0467_),
    .A(net761),
    .B(net757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2236_ (.Y(_0468_),
    .A(_0464_),
    .B(_0467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2237_ (.Y(_0469_),
    .A(net763),
    .B(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2238_ (.Y(_0470_),
    .A(_0456_),
    .B(_0469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2239_ (.Y(_0471_),
    .A(_0468_),
    .B(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2240_ (.Y(_0472_),
    .A(\u_usb_cdc.u_sie.data_q[5] ),
    .B(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2241_ (.Y(_0473_),
    .B1(_0471_),
    .B2(_0472_),
    .A2(_0466_),
    .A1(_1960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2242_ (.A0(_0471_),
    .A1(_0472_),
    .S(\u_usb_cdc.u_sie.data_q[7] ),
    .X(_0474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2243_ (.Y(_0475_),
    .A(\u_usb_cdc.u_sie.data_q[4] ),
    .B(_0468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2244_ (.Y(_0476_),
    .A(_0466_),
    .B(_0475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2245_ (.B1(_0476_),
    .VDD(VPWR),
    .Y(_0477_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_sie.data_q[6] ),
    .A2(_0475_));
 sg13g2_and4_1 _2246_ (.A(_0463_),
    .B(_0473_),
    .C(_0474_),
    .D(_0477_),
    .X(_0478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2247_ (.A(_0455_),
    .B(_0478_),
    .X(_0479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2248_ (.Y(_0480_),
    .B(_0479_),
    .A_N(_0453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2249_ (.Y(_0481_),
    .B(_0478_),
    .A_N(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2250_ (.Y(_0482_),
    .B(_0480_),
    .A_N(_0441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2251_ (.B(net766),
    .A(\u_usb_cdc.u_sie.crc16_q[14] ),
    .X(_0483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2252_ (.B(net767),
    .A(\u_usb_cdc.u_sie.crc16_q[15] ),
    .X(_0484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2253_ (.Y(_0485_),
    .A(_0483_),
    .B(_0484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2254_ (.Y(_0486_),
    .A(net920),
    .B(\u_usb_cdc.u_sie.data_q[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2255_ (.B(\u_usb_cdc.u_sie.data_q[3] ),
    .A(net913),
    .X(_0487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2256_ (.Y(_0488_),
    .A(_0486_),
    .B(_0487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2257_ (.B(_0487_),
    .A(_0486_),
    .X(_0489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2258_ (.Y(_0490_),
    .A(_0485_),
    .B(_0488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2259_ (.Y(_0491_),
    .A(\u_usb_cdc.u_sie.crc16_q[13] ),
    .B(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2260_ (.Y(_0492_),
    .A(net888),
    .B(\u_usb_cdc.u_sie.data_q[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2261_ (.Y(_0493_),
    .A(net967),
    .B(\u_usb_cdc.u_sie.data_q[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2262_ (.Y(_0494_),
    .A(_0492_),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2263_ (.B(_0494_),
    .A(_0491_),
    .X(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2264_ (.B(_0491_),
    .A(_0487_),
    .X(_0496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2265_ (.Y(_0497_),
    .A(_0490_),
    .B(_0495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2266_ (.Y(_0498_),
    .A(_1962_),
    .B(_0485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2267_ (.Y(_0499_),
    .A(\u_usb_cdc.u_sie.crc16_q[1] ),
    .B(_0484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2268_ (.B(_0491_),
    .A(_0483_),
    .X(_0500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2269_ (.Y(_0501_),
    .A(net915),
    .B(\u_usb_cdc.u_sie.data_q[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2270_ (.A(_0501_),
    .B_N(_0492_),
    .Y(_0502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2271_ (.A(\u_usb_cdc.u_sie.crc16_q[3] ),
    .B(\u_usb_cdc.u_sie.crc16_q[2] ),
    .Y(_0503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2272_ (.A(\u_usb_cdc.u_sie.crc16_q[5] ),
    .B(\u_usb_cdc.u_sie.crc16_q[4] ),
    .C(\u_usb_cdc.u_sie.crc16_q[7] ),
    .D(\u_usb_cdc.u_sie.crc16_q[6] ),
    .Y(_0504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2273_ (.Y(_0505_),
    .A(_0486_),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2274_ (.Y(_0506_),
    .B(net840),
    .A_N(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2275_ (.B(_0500_),
    .C(_0505_),
    .A(_0499_),
    .Y(_0507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2276_ (.B(_0502_),
    .C(_0503_),
    .A(_0496_),
    .Y(_0508_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0504_));
 sg13g2_nor4_1 _2277_ (.A(_0488_),
    .B(_0494_),
    .C(_0507_),
    .D(_0508_),
    .Y(_0509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2278_ (.B(_0498_),
    .C(_0509_),
    .A(_0497_),
    .Y(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2279_ (.VDD(VPWR),
    .Y(_0511_),
    .A(_0510_),
    .VSS(VGND));
 sg13g2_nand2_1 _2280_ (.Y(_0512_),
    .A(net841),
    .B(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2281_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0513_),
    .B(_0512_),
    .A(net750));
 sg13g2_nor2_1 _2282_ (.A(net768),
    .B(\u_usb_cdc.endp[1] ),
    .Y(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2283_ (.A(net769),
    .B_N(_2015_),
    .Y(_0515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2284_ (.Y(_0516_),
    .B(net710),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net768));
 sg13g2_nand2_1 _2285_ (.Y(_0517_),
    .A(\u_usb_cdc.ctrl_stall ),
    .B(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2286_ (.B(\u_usb_cdc.ctrl_stall ),
    .C(net640),
    .A(net847),
    .Y(_0518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2287_ (.A(\u_usb_cdc.u_sie.phy_state_q[2] ),
    .B(\u_usb_cdc.u_sie.phy_state_q[5] ),
    .C(\u_usb_cdc.u_sie.phy_state_q[3] ),
    .Y(_0519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2288_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0050_),
    .A2(_0519_),
    .Y(_0520_),
    .B1(net751));
 sg13g2_nor2_1 _2289_ (.A(net753),
    .B(net599),
    .Y(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2290_ (.A(net750),
    .B(net752),
    .C(net596),
    .Y(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2291_ (.Y(_0523_),
    .A(net844),
    .B(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2292_ (.B(net779),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .X(_0524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2293_ (.B(net787),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .X(_0525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2294_ (.B(net772),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .X(_0526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2295_ (.B(\u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .A(net778),
    .X(_0527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2296_ (.B(net793),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .X(_0528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2297_ (.B(net775),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .X(_0529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2298_ (.B(net790),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .X(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2299_ (.A(_0524_),
    .B(_0528_),
    .C(_0529_),
    .Y(_0531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2300_ (.A(_0525_),
    .B(_0526_),
    .C(_0527_),
    .D(_0530_),
    .Y(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2301_ (.Y(_0533_),
    .B(net788),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net785));
 sg13g2_nand2b_1 _2302_ (.Y(_0534_),
    .B(net788),
    .A_N(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2303_ (.A(net791),
    .B(net787),
    .C(net779),
    .Y(_0535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2304_ (.A(net790),
    .B(_0535_),
    .X(_0536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2305_ (.Y(_0537_),
    .B(net776),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net775));
 sg13g2_nor3_1 _2306_ (.A(net772),
    .B(_1926_),
    .C(_0537_),
    .Y(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2307_ (.Y(_0539_),
    .B(net791),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net784));
 sg13g2_and2_1 _2308_ (.A(net793),
    .B(net789),
    .X(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2309_ (.Y(_0541_),
    .A(net791),
    .B(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2310_ (.A(net784),
    .B(_0541_),
    .Y(_0542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2311_ (.B(net788),
    .C(net791),
    .Y(_0543_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net784));
 sg13g2_nor2_1 _2312_ (.A(net780),
    .B(_0543_),
    .Y(_0544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2313_ (.A(net776),
    .B(net773),
    .Y(_0545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2314_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0546_),
    .B(net775),
    .A(net776));
 sg13g2_nand2_1 _2315_ (.Y(_0547_),
    .A(net772),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2316_ (.A(net779),
    .B(_0543_),
    .C(_0546_),
    .D(_0547_),
    .Y(_0548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2317_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0538_),
    .C1(_0548_),
    .B1(_0536_),
    .A1(_0531_),
    .Y(_0549_),
    .A2(_0532_));
 sg13g2_nand2b_1 _2318_ (.Y(_0550_),
    .B(net541),
    .A_N(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _2319_ (.A(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .B(\u_usb_cdc.ctrl_stall ),
    .C(\u_usb_cdc.u_ctrl_endp.state_q[5] ),
    .D(_0550_),
    .X(_0551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2320_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0552_),
    .B(net850),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[1] ));
 sg13g2_nor2b_1 _2321_ (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .B_N(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .Y(_0553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2322_ (.A(net849),
    .B(_0551_),
    .C(_0552_),
    .D(_0553_),
    .Y(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2323_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0555_),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .A(net769));
 sg13g2_a21oi_2 _2324_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0555_),
    .Y(_0556_),
    .A2(_0554_),
    .A1(_0549_));
 sg13g2_nand2b_1 _2325_ (.Y(_0557_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2326_ (.Y(_0558_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ),
    .A_N(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2327_ (.Y(_0559_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ),
    .B(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2328_ (.Y(_0560_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2329_ (.B(_0558_),
    .C(_0560_),
    .A(\u_usb_cdc.endp[0] ),
    .Y(_0561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2330_ (.Y(_0562_),
    .B1(_1924_),
    .B2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ),
    .A2(net809),
    .A1(_1922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2331_ (.B(_0559_),
    .C(_0562_),
    .A(_0557_),
    .Y(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2332_ (.B1(net710),
    .VDD(VPWR),
    .Y(_0564_),
    .VSS(VGND),
    .A1(_0561_),
    .A2(_0563_));
 sg13g2_nor2_1 _2333_ (.A(_0556_),
    .B(_0564_),
    .Y(_0565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2334_ (.A(\u_usb_cdc.endp[1] ),
    .B_N(net768),
    .Y(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2335_ (.A(net769),
    .B(_2015_),
    .X(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2336_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net84),
    .C1(_0565_),
    .B1(net638),
    .A1(net164),
    .Y(_0568_),
    .A2(net640));
 sg13g2_nand2_1 _2337_ (.Y(_0569_),
    .A(net847),
    .B(_0517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2338_ (.A(_2017_),
    .B(_0569_),
    .Y(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2339_ (.A(net594),
    .B(_0570_),
    .X(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2340_ (.Y(_0572_),
    .A(net594),
    .B(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2341_ (.Y(_0573_),
    .A(_0568_),
    .B(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2342_ (.B1(_0573_),
    .VDD(VPWR),
    .Y(_0574_),
    .VSS(VGND),
    .A1(net141),
    .A2(net601));
 sg13g2_a21oi_1 _2343_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net847),
    .A2(_2017_),
    .Y(_0575_),
    .B1(_0520_));
 sg13g2_and2_1 _2344_ (.A(_0513_),
    .B(_0575_),
    .X(_0576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2345_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0482_),
    .A2(_0576_),
    .Y(_0577_),
    .B1(net752));
 sg13g2_or2_1 _2346_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0578_),
    .B(_0510_),
    .A(_0506_));
 sg13g2_nor2_1 _2347_ (.A(net710),
    .B(_0578_),
    .Y(_0579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2348_ (.A(net836),
    .B(net837),
    .C(_0577_),
    .D(_0579_),
    .Y(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2349_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0518_),
    .A2(net987),
    .Y(_0581_),
    .B1(net596));
 sg13g2_a22oi_1 _2350_ (.Y(_0582_),
    .B1(net844),
    .B2(_0522_),
    .A2(net745),
    .A1(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2351_ (.VDD(VPWR),
    .Y(_0583_),
    .A(_0582_),
    .VSS(VGND));
 sg13g2_nor3_1 _2352_ (.A(_0574_),
    .B(net988),
    .C(_0583_),
    .Y(_0063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2353_ (.B(net327),
    .C(net321),
    .A(net376),
    .Y(_0584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2354_ (.A(\u_usb_cdc.u_sie.in_byte_q[3] ),
    .B(_2017_),
    .C(_0584_),
    .Y(_0585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2355_ (.A(_1919_),
    .B(_0585_),
    .Y(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2356_ (.A(_1919_),
    .B(_0556_),
    .C(_0564_),
    .D(_0585_),
    .Y(_0587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2357_ (.A(net850),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .C(_0551_),
    .X(_0588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2358_ (.A(_0516_),
    .B(_0588_),
    .Y(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2359_ (.Y(_0590_),
    .B(_0565_),
    .A_N(_0589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2360_ (.A(_0556_),
    .B(_0564_),
    .C(_0569_),
    .D(_0589_),
    .Y(_0591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2361_ (.B1(_0435_),
    .VDD(VPWR),
    .Y(_0592_),
    .VSS(VGND),
    .A1(_0587_),
    .A2(_0591_));
 sg13g2_nor2_1 _2362_ (.A(\u_usb_cdc.sie_in_data_ack ),
    .B(\u_usb_cdc.sie_in_req ),
    .Y(_0593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2363_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0592_),
    .A2(_0593_),
    .Y(_0594_),
    .B1(_0516_));
 sg13g2_nand2_2 _2364_ (.Y(_0595_),
    .A(\u_usb_cdc.sie_in_req ),
    .B(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2365_ (.B1(_0595_),
    .VDD(VPWR),
    .Y(_0596_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .A2(\u_usb_cdc.u_ctrl_endp.state_q[5] ));
 sg13g2_a21oi_1 _2366_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1918_),
    .A2(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .Y(_0597_),
    .B1(\u_usb_cdc.u_ctrl_endp.state_q[2] ));
 sg13g2_a221oi_1 _2367_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0597_),
    .C1(_0516_),
    .B1(_0596_),
    .A1(_0592_),
    .Y(_0598_),
    .A2(_0593_));
 sg13g2_nand2b_1 _2368_ (.Y(_0599_),
    .B(net750),
    .A_N(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2369_ (.Y(_0600_),
    .A(net751),
    .B(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2370_ (.A(net752),
    .B(_0600_),
    .Y(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2371_ (.A(_0601_),
    .Y(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2372_ (.B(net430),
    .C(net354),
    .A(net156),
    .Y(_0603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2373_ (.A(net755),
    .B(_0601_),
    .Y(_0604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2374_ (.Y(_0605_),
    .B1(_0604_),
    .B2(_1931_),
    .A2(_0603_),
    .A1(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2375_ (.A(net640),
    .B(_0605_),
    .X(_0606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2376_ (.A(net849),
    .B(net471),
    .C(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .Y(_0607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2377_ (.B1(_0607_),
    .VDD(VPWR),
    .Y(_0608_),
    .VSS(VGND),
    .A1(_1928_),
    .A2(_0602_));
 sg13g2_nand2_1 _2378_ (.Y(_0609_),
    .A(_0606_),
    .B(_0608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2379_ (.A(_0598_),
    .B_N(_0609_),
    .Y(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2380_ (.Y(_0611_),
    .B(_0609_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0598_));
 sg13g2_nand2_2 _2381_ (.Y(_0612_),
    .A(net755),
    .B(_0606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2382_ (.B(\u_usb_cdc.u_sie.pid_q[3] ),
    .C(_0451_),
    .A(net1053),
    .Y(_0613_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0606_));
 sg13g2_and2_1 _2383_ (.A(_0612_),
    .B(_0613_),
    .X(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2384_ (.Y(_0615_),
    .A(_0612_),
    .B(_0613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2385_ (.B1(_0614_),
    .VDD(VPWR),
    .Y(_0616_),
    .VSS(VGND),
    .A1(_0594_),
    .A2(_0606_));
 sg13g2_nor2_2 _2386_ (.A(_0611_),
    .B(_0616_),
    .Y(_0617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2387_ (.B1(net743),
    .VDD(VPWR),
    .Y(_0618_),
    .VSS(VGND),
    .A1(_0594_),
    .A2(_0606_));
 sg13g2_inv_2 _2388_ (.Y(_0619_),
    .A(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2389_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0620_),
    .B(net590),
    .A(_0615_));
 sg13g2_nand3b_1 _2390_ (.B(_0609_),
    .C(_0614_),
    .Y(_0621_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0598_));
 sg13g2_nor2_1 _2391_ (.A(net590),
    .B(_0621_),
    .Y(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2392_ (.Y(_0623_),
    .A(net743),
    .B(_0617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2393_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_usb_cdc.sie_in_req ),
    .A2(net640),
    .Y(_0624_),
    .B1(\u_usb_cdc.sie_in_data_ack ));
 sg13g2_nand2_1 _2394_ (.Y(_0625_),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .B(_0624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2395_ (.B(net541),
    .C(_0625_),
    .Y(_0626_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net849));
 sg13g2_nor2_1 _2396_ (.A(_0550_),
    .B(_0552_),
    .Y(_0627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2397_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0607_),
    .A2(_0627_),
    .Y(_0628_),
    .B1(_0612_));
 sg13g2_nor2_1 _2398_ (.A(net541),
    .B(_0619_),
    .Y(_0629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2399_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net742),
    .C1(_0629_),
    .B1(_0628_),
    .A1(net589),
    .Y(_0062_),
    .A2(_0626_));
 sg13g2_nand2_2 _2400_ (.Y(_0630_),
    .A(net850),
    .B(_0601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2401_ (.A(_0611_),
    .B(_0616_),
    .C(net624),
    .Y(_0631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2402_ (.B(_0601_),
    .C(_0617_),
    .A(net968),
    .Y(_0632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2403_ (.A(net772),
    .B(_0546_),
    .Y(_0633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2404_ (.A(net779),
    .B(net772),
    .C(_0546_),
    .Y(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2405_ (.Y(_0635_),
    .B(_0633_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net779));
 sg13g2_nand3_1 _2406_ (.B(_0542_),
    .C(_0634_),
    .A(net744),
    .Y(_0636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2407_ (.A(_0611_),
    .B(_0616_),
    .C(net624),
    .Y(_0637_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0636_));
 sg13g2_and2_1 _2408_ (.A(_0536_),
    .B(_0633_),
    .X(_0638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2409_ (.Y(_0639_),
    .A(_0536_),
    .B(_0633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2410_ (.Y(_0640_),
    .A(net743),
    .B(_0638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2411_ (.A(_0611_),
    .B(_0616_),
    .C(_0630_),
    .Y(_0641_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0640_));
 sg13g2_nor2_1 _2412_ (.A(_0637_),
    .B(_0641_),
    .Y(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2413_ (.A(net849),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .C(_0551_),
    .Y(_0643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2414_ (.VDD(VPWR),
    .Y(_0644_),
    .A(_0643_),
    .VSS(VGND));
 sg13g2_nand2_2 _2415_ (.Y(_0645_),
    .A(net787),
    .B(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2416_ (.VDD(VPWR),
    .Y(_0646_),
    .A(_0645_),
    .VSS(VGND));
 sg13g2_nor2b_2 _2417_ (.A(net782),
    .B_N(net784),
    .Y(_0647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2418_ (.A(_0534_),
    .B(_0645_),
    .Y(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2419_ (.Y(_0649_),
    .A(net743),
    .B(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _2420_ (.A(_0611_),
    .B(_0616_),
    .C(_0630_),
    .D(_0649_),
    .X(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2421_ (.X(_0651_),
    .A(net588),
    .B(_0643_),
    .C(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2422_ (.Y(_0652_),
    .A(net792),
    .B(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2423_ (.A2(_0540_),
    .A1(net785),
    .B1(net781),
    .X(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2424_ (.A(net777),
    .B(_0653_),
    .Y(_0654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2425_ (.Y(_0655_),
    .A(net785),
    .B(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2426_ (.B1(net776),
    .VDD(VPWR),
    .Y(_0656_),
    .VSS(VGND),
    .A1(_0534_),
    .A2(_0655_));
 sg13g2_nand2b_2 _2427_ (.Y(_0657_),
    .B(net780),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net777));
 sg13g2_nor2b_1 _2428_ (.A(net774),
    .B_N(net781),
    .Y(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2429_ (.B1(_0656_),
    .VDD(VPWR),
    .Y(_0659_),
    .VSS(VGND),
    .A1(_0542_),
    .A2(_0657_));
 sg13g2_nor3_1 _2430_ (.A(_0654_),
    .B(_0658_),
    .C(_0659_),
    .Y(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2431_ (.Y(_0661_),
    .A(_0633_),
    .B(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2432_ (.A(net590),
    .B(_0621_),
    .C(net624),
    .Y(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2433_ (.A(net590),
    .B(_0621_),
    .C(net624),
    .D(_0661_),
    .Y(_0663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2434_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0635_),
    .A2(_0662_),
    .Y(_0664_),
    .B1(_0663_));
 sg13g2_nor2b_2 _2435_ (.A(_0601_),
    .B_N(net850),
    .Y(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2436_ (.Y(_0666_),
    .A(net850),
    .B(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2437_ (.A(net590),
    .B(_0621_),
    .C(_0666_),
    .Y(_0667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2438_ (.A(net791),
    .B(net790),
    .Y(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2439_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0669_),
    .B(net788),
    .A(net791));
 sg13g2_nand2_1 _2440_ (.Y(_0670_),
    .A(_1925_),
    .B(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2441_ (.A(_0645_),
    .B(_0669_),
    .Y(_0671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2442_ (.Y(_0672_),
    .A(_0646_),
    .B(_0668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2443_ (.A(net590),
    .B(_0621_),
    .C(net624),
    .Y(_0673_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0672_));
 sg13g2_nor2b_1 _2444_ (.A(net788),
    .B_N(net791),
    .Y(_0674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2445_ (.Y(_0675_),
    .A(net791),
    .B(_1925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2446_ (.A(_0645_),
    .B(_0675_),
    .Y(_0676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2447_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0662_),
    .C1(_0673_),
    .B1(_0676_),
    .A1(net588),
    .Y(_0677_),
    .A2(_0665_));
 sg13g2_nand3_1 _2448_ (.B(_0664_),
    .C(_0677_),
    .A(_0651_),
    .Y(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2449_ (.B(_0651_),
    .C(_0664_),
    .A(_0642_),
    .Y(_0679_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0677_));
 sg13g2_a221oi_1 _2450_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0644_),
    .C1(net590),
    .B1(net588),
    .A1(net756),
    .Y(_0680_),
    .A2(_0606_));
 sg13g2_a221oi_1 _2451_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0613_),
    .C1(net591),
    .B1(_0610_),
    .A1(net756),
    .Y(_0681_),
    .A2(_0606_));
 sg13g2_nor2_2 _2452_ (.A(net760),
    .B(net761),
    .Y(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2453_ (.B1(_0682_),
    .VDD(VPWR),
    .Y(_0683_),
    .VSS(VGND),
    .A1(net723),
    .A2(net721));
 sg13g2_nor3_1 _2454_ (.A(net759),
    .B(net758),
    .C(_0683_),
    .Y(_0684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2455_ (.A(net787),
    .B(_0669_),
    .Y(_0685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2456_ (.Y(_0686_),
    .A(_0634_),
    .B(_0685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2457_ (.A(net759),
    .B(net758),
    .C(_0683_),
    .D(_0686_),
    .Y(_0687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2458_ (.Y(_0061_),
    .B1(_0687_),
    .B2(_0662_),
    .A2(_0679_),
    .A1(_2005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2459_ (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .B(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .X(\u_usb_cdc.configured_o ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2460_ (.A(net298),
    .B(net757),
    .C(\u_usb_cdc.sie_out_data[6] ),
    .Y(_0688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2461_ (.A(_1914_),
    .B(_0688_),
    .X(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2462_ (.A(_1913_),
    .B(_0689_),
    .X(_0690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2463_ (.Y(_0691_),
    .A(_0682_),
    .B(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2464_ (.A(net762),
    .B(_0691_),
    .Y(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2465_ (.B(_0682_),
    .C(_0689_),
    .A(net721),
    .Y(_0693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2466_ (.A(net723),
    .B(_0693_),
    .Y(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2467_ (.Y(_0695_),
    .A(net763),
    .B(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2468_ (.B1(_0680_),
    .VDD(VPWR),
    .Y(_0696_),
    .VSS(VGND),
    .A1(_0650_),
    .A2(_0695_));
 sg13g2_nor2_1 _2469_ (.A(net763),
    .B(_0693_),
    .Y(_0697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2470_ (.Y(_0698_),
    .A(net723),
    .B(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2471_ (.B(_0646_),
    .C(_0662_),
    .A(_1925_),
    .Y(_0699_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net622));
 sg13g2_nand2_1 _2472_ (.Y(_0700_),
    .A(_0637_),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2473_ (.B1(net623),
    .VDD(VPWR),
    .Y(_0701_),
    .VSS(VGND),
    .A1(_0637_),
    .A2(_0641_));
 sg13g2_nand2_1 _2474_ (.Y(_0702_),
    .A(_0663_),
    .B(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2475_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net588),
    .C1(_0681_),
    .B1(_0665_),
    .A1(_0635_),
    .Y(_0703_),
    .A2(_0662_));
 sg13g2_nand4_1 _2476_ (.B(_0701_),
    .C(_0702_),
    .A(_0699_),
    .Y(_0704_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0703_));
 sg13g2_o21ai_1 _2477_ (.B1(net874),
    .VDD(VPWR),
    .Y(_0705_),
    .VSS(VGND),
    .A1(_0696_),
    .A2(_0704_));
 sg13g2_nand2b_2 _2478_ (.Y(_0706_),
    .B(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net413));
 sg13g2_nand2_1 _2479_ (.Y(_0707_),
    .A(\u_usb_cdc.sie_out_data[3] ),
    .B(_0690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2480_ (.B(_0690_),
    .C(_0706_),
    .A(\u_usb_cdc.sie_out_data[3] ),
    .Y(_0708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2481_ (.A(net880),
    .B(net953),
    .Y(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2482_ (.Y(_0710_),
    .A(net794),
    .B(_0709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _2483_ (.A(net763),
    .B(net762),
    .C(_0708_),
    .D(_0710_),
    .X(_0711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2484_ (.B(_0610_),
    .C(_0613_),
    .A(net850),
    .Y(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2485_ (.A(net752),
    .B(net756),
    .Y(_0713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2486_ (.A(net756),
    .B(_0602_),
    .Y(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2487_ (.Y(_0715_),
    .A(net641),
    .B(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _2488_ (.A(net492),
    .B(_0712_),
    .C(_0715_),
    .X(_0716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2489_ (.A(net938),
    .B(_0716_),
    .Y(_0717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2490_ (.A(net789),
    .B(_0539_),
    .Y(_0718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2491_ (.A(net787),
    .B(net715),
    .C(_0635_),
    .Y(_0719_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0675_));
 sg13g2_nand2_2 _2492_ (.Y(_0720_),
    .A(_0717_),
    .B(_0719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2493_ (.B1(_0705_),
    .VDD(VPWR),
    .Y(_0005_),
    .VSS(VGND),
    .A1(_0711_),
    .A2(_0720_));
 sg13g2_nand2_1 _2494_ (.Y(_0721_),
    .A(net942),
    .B(_0679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2495_ (.B(\u_usb_cdc.sie_out_data[2] ),
    .C(_0689_),
    .A(net720),
    .Y(_0722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2496_ (.Y(_0723_),
    .A(_0707_),
    .B(_0722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2497_ (.Y(_0724_),
    .B(_0723_),
    .A_N(_0459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2498_ (.X(_0725_),
    .A(_0693_),
    .B(_0711_),
    .C(_0724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2499_ (.Y(_0726_),
    .A(net794),
    .B(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2500_ (.Y(_0727_),
    .A(net723),
    .B(\u_usb_cdc.sie_out_data[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2501_ (.A(_0707_),
    .B(_0727_),
    .Y(_0728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2502_ (.B(_1937_),
    .C(net794),
    .A(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .Y(_0729_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\u_usb_cdc.configured_o ));
 sg13g2_a22oi_1 _2503_ (.Y(_0730_),
    .B1(_0728_),
    .B2(_0729_),
    .A2(_0726_),
    .A1(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2504_ (.Y(_0731_),
    .B(_0730_),
    .A_N(_0725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2505_ (.Y(_0732_),
    .A(_1938_),
    .B(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2506_ (.B1(_0709_),
    .VDD(VPWR),
    .Y(_0733_),
    .VSS(VGND),
    .A1(_1938_),
    .A2(_0722_));
 sg13g2_nor3_1 _2507_ (.A(net880),
    .B(net953),
    .C(net794),
    .Y(_0734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2508_ (.Y(_0735_),
    .B1(_0733_),
    .B2(_0723_),
    .A2(_0732_),
    .A1(_0690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2509_ (.B(net721),
    .C(_0719_),
    .A(net764),
    .Y(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2510_ (.VDD(VPWR),
    .Y(_0737_),
    .A(_0736_),
    .VSS(VGND));
 sg13g2_nor2_1 _2511_ (.A(_0735_),
    .B(_0736_),
    .Y(_0738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2512_ (.A(_0722_),
    .B(_0727_),
    .Y(_0739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2513_ (.A(_0719_),
    .B(_0739_),
    .X(_0740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2514_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0710_),
    .C1(_0738_),
    .B1(_0740_),
    .A1(_0719_),
    .Y(_0741_),
    .A2(_0731_));
 sg13g2_nor2_1 _2515_ (.A(_0716_),
    .B(_0741_),
    .Y(_0742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2516_ (.B(net851),
    .C(_0638_),
    .A(net743),
    .Y(_0743_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0693_));
 sg13g2_nor2_1 _2517_ (.A(_1942_),
    .B(_0636_),
    .Y(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2518_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0745_),
    .B(_0727_),
    .A(_0691_));
 sg13g2_nand3_1 _2519_ (.B(_0744_),
    .C(_0745_),
    .A(_0695_),
    .Y(_0746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2520_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .B(net851),
    .Y(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2521_ (.Y(_0748_),
    .A(_1941_),
    .B(_0747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2522_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0749_),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[4] ));
 sg13g2_nor3_1 _2523_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .B(_0748_),
    .C(_0749_),
    .Y(_0750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2524_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .Y(_0751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2525_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .C(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .Y(_0752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2526_ (.B(_0751_),
    .C(_0752_),
    .A(_0750_),
    .Y(_0753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2527_ (.A(_0649_),
    .B(net622),
    .C(_0749_),
    .Y(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2528_ (.Y(_0755_),
    .B1(_0754_),
    .B2(_0748_),
    .A2(_0753_),
    .A1(_0719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2529_ (.B(_0746_),
    .C(_0755_),
    .A(_0743_),
    .Y(_0756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2530_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0631_),
    .A2(_0756_),
    .Y(_0757_),
    .B1(_0742_));
 sg13g2_nand4_1 _2531_ (.B(_0682_),
    .C(\u_usb_cdc.configured_o ),
    .A(\u_usb_cdc.sie_out_data[5] ),
    .Y(_0758_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0688_));
 sg13g2_nand4_1 _2532_ (.B(net641),
    .C(_0714_),
    .A(net492),
    .Y(_0759_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0719_));
 sg13g2_nor2_1 _2533_ (.A(_0712_),
    .B(_0759_),
    .Y(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2534_ (.Y(_0761_),
    .A(net787),
    .B(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2535_ (.B1(_0761_),
    .VDD(VPWR),
    .Y(_0762_),
    .VSS(VGND),
    .A1(net784),
    .A2(_0540_));
 sg13g2_or2_1 _2536_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0763_),
    .B(_0762_),
    .A(_0635_));
 sg13g2_a21oi_1 _2537_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0661_),
    .A2(_0763_),
    .Y(_0764_),
    .B1(_0750_));
 sg13g2_or3_1 _2538_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .B(net851),
    .C(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .X(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2539_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0671_),
    .A2(_0765_),
    .Y(_0766_),
    .B1(_0764_));
 sg13g2_nand2_1 _2540_ (.Y(_0767_),
    .A(_1936_),
    .B(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2541_ (.A(net721),
    .B(net757),
    .Y(_0768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2542_ (.A(_0683_),
    .B(_0767_),
    .C(_0768_),
    .Y(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2543_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net764),
    .A2(_1936_),
    .Y(_0770_),
    .B1(\u_usb_cdc.u_ctrl_endp.rec_q[1] ));
 sg13g2_a21oi_1 _2544_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0692_),
    .A2(_0770_),
    .Y(_0771_),
    .B1(_0769_));
 sg13g2_nor2b_1 _2545_ (.A(_0769_),
    .B_N(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .Y(_0772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2546_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .C1(_0772_),
    .B1(_0771_),
    .A1(\u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .Y(_0773_),
    .A2(_0693_));
 sg13g2_nor2_1 _2547_ (.A(_0672_),
    .B(_0773_),
    .Y(_0774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2548_ (.Y(_0775_),
    .B1(_0749_),
    .B2(_0695_),
    .A2(_0745_),
    .A1(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2549_ (.A(_0775_),
    .B_N(_0648_),
    .Y(_0776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2550_ (.B1(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .VDD(VPWR),
    .Y(_0777_),
    .VSS(VGND),
    .A1(_0698_),
    .A2(_0767_));
 sg13g2_or3_1 _2551_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .C(_0749_),
    .X(_0778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2552_ (.Y(_0779_),
    .B1(_0698_),
    .B2(_0778_),
    .A2(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .A1(net757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2553_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0777_),
    .A2(_0779_),
    .Y(_0780_),
    .B1(_0639_));
 sg13g2_or4_1 _2554_ (.A(net790),
    .B(_0645_),
    .C(net622),
    .D(_0751_),
    .X(_0781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2555_ (.B1(_0781_),
    .VDD(VPWR),
    .Y(_0782_),
    .VSS(VGND),
    .A1(_0684_),
    .A2(_0686_));
 sg13g2_nor4_1 _2556_ (.A(_0774_),
    .B(_0776_),
    .C(_0780_),
    .D(_0782_),
    .Y(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2557_ (.B1(_0783_),
    .VDD(VPWR),
    .Y(_0784_),
    .VSS(VGND),
    .A1(net622),
    .A2(_0766_));
 sg13g2_a22oi_1 _2558_ (.Y(_0785_),
    .B1(_0784_),
    .B2(_0662_),
    .A2(_0760_),
    .A1(_0758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2559_ (.B(_0757_),
    .C(_0785_),
    .A(_0721_),
    .Y(_0004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2560_ (.Y(_0786_),
    .A(_0641_),
    .B(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2561_ (.A(_0649_),
    .B(_0698_),
    .C(_0749_),
    .Y(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2562_ (.Y(_0788_),
    .A(_0631_),
    .B(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2563_ (.B(_0786_),
    .C(_0788_),
    .A(_0680_),
    .Y(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2564_ (.B1(net513),
    .VDD(VPWR),
    .Y(_0790_),
    .VSS(VGND),
    .A1(_0704_),
    .A2(_0789_));
 sg13g2_nand3_1 _2565_ (.B(_0734_),
    .C(_0737_),
    .A(_0717_),
    .Y(_0791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2566_ (.B1(_0790_),
    .VDD(VPWR),
    .Y(_0006_),
    .VSS(VGND),
    .A1(_0708_),
    .A2(_0791_));
 sg13g2_nor3_1 _2567_ (.A(_0610_),
    .B(_0615_),
    .C(net591),
    .Y(_0792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2568_ (.Y(_0793_),
    .A(_0643_),
    .B(_0666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2569_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net588),
    .C1(_0792_),
    .B1(_0793_),
    .A1(_0663_),
    .Y(_0794_),
    .A2(net622));
 sg13g2_nand3_1 _2570_ (.B(_0788_),
    .C(_0794_),
    .A(_0700_),
    .Y(_0795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2571_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0635_),
    .A2(_0662_),
    .Y(_0796_),
    .B1(_0620_));
 sg13g2_nand4_1 _2572_ (.B(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .C(_0641_),
    .A(_1936_),
    .Y(_0797_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net623));
 sg13g2_nand2_1 _2573_ (.Y(_0798_),
    .A(_0673_),
    .B(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2574_ (.B(_0676_),
    .C(net622),
    .A(_0662_),
    .Y(_0799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2575_ (.B(_0797_),
    .C(_0798_),
    .A(_0796_),
    .Y(_0800_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0799_));
 sg13g2_o21ai_1 _2576_ (.B1(net483),
    .VDD(VPWR),
    .Y(_0801_),
    .VSS(VGND),
    .A1(_0795_),
    .A2(_0800_));
 sg13g2_nand3b_1 _2577_ (.B(_0694_),
    .C(_0706_),
    .Y(_0802_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sg13g2_o21ai_1 _2578_ (.B1(_0801_),
    .VDD(VPWR),
    .Y(_0007_),
    .VSS(VGND),
    .A1(_0720_),
    .A2(_0802_));
 sg13g2_nand2_1 _2579_ (.Y(_0803_),
    .A(net719),
    .B(_0641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2580_ (.B(_0796_),
    .C(_0803_),
    .A(_0699_),
    .Y(_0804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2581_ (.B1(net957),
    .VDD(VPWR),
    .Y(_0805_),
    .VSS(VGND),
    .A1(_0795_),
    .A2(_0804_));
 sg13g2_o21ai_1 _2582_ (.B1(_0805_),
    .VDD(VPWR),
    .Y(_0008_),
    .VSS(VGND),
    .A1(_0722_),
    .A2(_0791_));
 sg13g2_nor3_1 _2583_ (.A(_0637_),
    .B(_0641_),
    .C(_0667_),
    .Y(_0806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2584_ (.B(_0664_),
    .C(_0699_),
    .A(_0651_),
    .Y(_0807_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0806_));
 sg13g2_nor4_1 _2585_ (.A(_1942_),
    .B(_0632_),
    .C(_0636_),
    .D(_0745_),
    .Y(_0808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2586_ (.A2(_0807_),
    .A1(net974),
    .B1(_0808_),
    .X(_0009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2587_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0641_),
    .A2(net622),
    .Y(_0809_),
    .B1(_0678_));
 sg13g2_nand4_1 _2588_ (.B(_0709_),
    .C(_0717_),
    .A(net794),
    .Y(_0810_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0740_));
 sg13g2_o21ai_1 _2589_ (.B1(_0810_),
    .VDD(VPWR),
    .Y(_0010_),
    .VSS(VGND),
    .A1(_1942_),
    .A2(_0809_));
 sg13g2_nor4_1 _2590_ (.A(_0048_),
    .B(_0712_),
    .C(_0758_),
    .D(_0759_),
    .Y(_0811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2591_ (.A2(_0679_),
    .A1(net411),
    .B1(_0811_),
    .X(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2592_ (.B(_0794_),
    .C(_0796_),
    .A(_0701_),
    .Y(_0812_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0799_));
 sg13g2_nand2_1 _2593_ (.Y(_0813_),
    .A(_0673_),
    .B(_0692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2594_ (.B1(_0813_),
    .VDD(VPWR),
    .Y(_0814_),
    .VSS(VGND),
    .A1(_0650_),
    .A2(_0695_));
 sg13g2_o21ai_1 _2595_ (.B1(net522),
    .VDD(VPWR),
    .Y(_0815_),
    .VSS(VGND),
    .A1(_0812_),
    .A2(_0814_));
 sg13g2_or3_1 _2596_ (.A(_0707_),
    .B(_0727_),
    .C(_0729_),
    .X(_0816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2597_ (.B1(_0815_),
    .VDD(VPWR),
    .Y(_0001_),
    .VSS(VGND),
    .A1(_0720_),
    .A2(_0816_));
 sg13g2_a21oi_1 _2598_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0595_),
    .A2(_0617_),
    .Y(_0817_),
    .B1(net591));
 sg13g2_nor3_1 _2599_ (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .B(\u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .C(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .Y(_0818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2600_ (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .B(\u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .C(\u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .D(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .Y(_0819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2601_ (.Y(_0820_),
    .A(_0818_),
    .B(_0819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2602_ (.Y(_0821_),
    .A(net779),
    .B(_0685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _2603_ (.A(net772),
    .B(net942),
    .C(_0546_),
    .D(_0821_),
    .X(_0822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2604_ (.VDD(VPWR),
    .Y(_0823_),
    .A(_0822_),
    .VSS(VGND));
 sg13g2_nor3_1 _2605_ (.A(net946),
    .B(_0666_),
    .C(_0822_),
    .Y(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2606_ (.Y(_0825_),
    .A(net588),
    .B(_0824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2607_ (.B(_0617_),
    .C(_0820_),
    .A(net742),
    .Y(_0826_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0824_));
 sg13g2_o21ai_1 _2608_ (.B1(_0826_),
    .VDD(VPWR),
    .Y(_0011_),
    .VSS(VGND),
    .A1(_1927_),
    .A2(_0817_));
 sg13g2_nand3b_1 _2609_ (.B(_0619_),
    .C(_0612_),
    .Y(_0827_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0613_));
 sg13g2_nand2_1 _2610_ (.Y(_0828_),
    .A(net968),
    .B(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2611_ (.B(_0827_),
    .C(_0828_),
    .A(_0632_),
    .Y(_0012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2612_ (.A(_1927_),
    .B(_0595_),
    .C(_0615_),
    .Y(_0829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2613_ (.B(_0610_),
    .C(_0829_),
    .A(net742),
    .Y(_0830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2614_ (.Y(_0831_),
    .B1(net589),
    .B2(net471),
    .A2(net591),
    .A1(net849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2615_ (.Y(_0013_),
    .A(_0830_),
    .B(_0831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2616_ (.Y(_0832_),
    .B1(_0827_),
    .B2(net1030),
    .A2(_0822_),
    .A1(_0667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2617_ (.Y(_0014_),
    .B(_0832_),
    .A_N(_0792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2618_ (.Y(_0833_),
    .A(net471),
    .B(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2619_ (.B1(_0833_),
    .VDD(VPWR),
    .Y(_0015_),
    .VSS(VGND),
    .A1(_0820_),
    .A2(_0825_));
 sg13g2_nor4_1 _2620_ (.A(\u_usb_cdc.sie_in_data_ack ),
    .B(_0549_),
    .C(_0595_),
    .D(_0615_),
    .Y(_0834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2621_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0610_),
    .C1(net591),
    .B1(_0834_),
    .A1(_0549_),
    .Y(_0835_),
    .A2(net589));
 sg13g2_nand4_1 _2622_ (.B(net588),
    .C(_0665_),
    .A(net946),
    .Y(_0836_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0823_));
 sg13g2_o21ai_1 _2623_ (.B1(net947),
    .VDD(VPWR),
    .Y(_0016_),
    .VSS(VGND),
    .A1(_1929_),
    .A2(_0835_));
 sg13g2_nor3_1 _2624_ (.A(_1918_),
    .B(_1929_),
    .C(_0549_),
    .Y(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2625_ (.A(_1928_),
    .B(_0624_),
    .Y(_0838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2626_ (.B1(net589),
    .VDD(VPWR),
    .Y(_0839_),
    .VSS(VGND),
    .A1(_0837_),
    .A2(_0838_));
 sg13g2_o21ai_1 _2627_ (.B1(_0839_),
    .VDD(VPWR),
    .Y(_0017_),
    .VSS(VGND),
    .A1(_1928_),
    .A2(_0619_));
 sg13g2_nand2_1 _2628_ (.Y(_0840_),
    .A(net847),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2629_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0841_),
    .B(_0481_),
    .A(_0453_));
 sg13g2_nand2_1 _2630_ (.Y(_0842_),
    .A(_0455_),
    .B(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2631_ (.B1(_0840_),
    .VDD(VPWR),
    .Y(_0020_),
    .VSS(VGND),
    .A1(_0841_),
    .A2(_0842_));
 sg13g2_nand2_1 _2632_ (.Y(_0843_),
    .A(net524),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2633_ (.Y(_0844_),
    .A(net750),
    .B(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2634_ (.B(net844),
    .C(net593),
    .A(net750),
    .Y(_0845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2635_ (.Y(_0846_),
    .A(\u_usb_cdc.addr[5] ),
    .B(\u_usb_cdc.u_sie.addr_q[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2636_ (.Y(_0847_),
    .A(\u_usb_cdc.addr[3] ),
    .B(\u_usb_cdc.u_sie.addr_q[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2637_ (.Y(_0848_),
    .A(\u_usb_cdc.addr[4] ),
    .B(\u_usb_cdc.u_sie.addr_q[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2638_ (.B(\u_usb_cdc.u_sie.addr_q[6] ),
    .A(\u_usb_cdc.addr[6] ),
    .X(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2639_ (.B(\u_usb_cdc.u_sie.addr_q[0] ),
    .A(\u_usb_cdc.addr[0] ),
    .X(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2640_ (.B(\u_usb_cdc.u_sie.addr_q[1] ),
    .A(\u_usb_cdc.addr[1] ),
    .X(_0851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2641_ (.B(\u_usb_cdc.u_sie.addr_q[2] ),
    .A(\u_usb_cdc.addr[2] ),
    .X(_0852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2642_ (.A(_0849_),
    .B(_0850_),
    .C(_0851_),
    .D(_0852_),
    .Y(_0853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2643_ (.B(_0847_),
    .C(_0848_),
    .A(_0846_),
    .Y(_0854_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0853_));
 sg13g2_o21ai_1 _2644_ (.B1(_0451_),
    .VDD(VPWR),
    .Y(_0855_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_sie.pid_q[2] ),
    .A2(_1935_));
 sg13g2_nor3_1 _2645_ (.A(net765),
    .B(_0454_),
    .C(_0855_),
    .Y(_0856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2646_ (.Y(_0857_),
    .A(net710),
    .B(_0856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2647_ (.Y(_0858_),
    .A(net767),
    .B(\u_usb_cdc.u_sie.data_q[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2648_ (.Y(_0859_),
    .A(net766),
    .B(\u_usb_cdc.u_sie.data_q[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2649_ (.Y(_0860_),
    .A(\u_usb_cdc.u_sie.data_q[3] ),
    .B(\u_usb_cdc.u_sie.data_q[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2650_ (.Y(_0861_),
    .A(net765),
    .B(\u_usb_cdc.u_sie.data_q[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _2651_ (.A(_0858_),
    .B(_0859_),
    .C(_0860_),
    .Y(_0862_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0861_));
 sg13g2_nand2_1 _2652_ (.Y(_0863_),
    .A(net767),
    .B(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2653_ (.A(_0854_),
    .B(_0857_),
    .C(_0863_),
    .Y(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2654_ (.Y(_0865_),
    .A(net766),
    .B(_0864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2655_ (.B1(_0843_),
    .VDD(VPWR),
    .Y(_0021_),
    .VSS(VGND),
    .A1(_0845_),
    .A2(_0865_));
 sg13g2_or3_1 _2656_ (.A(net766),
    .B(_0845_),
    .C(_0863_),
    .X(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2657_ (.B1(net561),
    .VDD(VPWR),
    .Y(_0022_),
    .VSS(VGND),
    .A1(_1974_),
    .A2(net601));
 sg13g2_nand2_2 _2658_ (.Y(_0867_),
    .A(net843),
    .B(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2659_ (.A(_0568_),
    .B_N(_0590_),
    .Y(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2660_ (.Y(_0869_),
    .B1(_0571_),
    .B2(_0868_),
    .A2(net596),
    .A1(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2661_ (.B1(_0869_),
    .VDD(VPWR),
    .Y(_0023_),
    .VSS(VGND),
    .A1(_0587_),
    .A2(_0867_));
 sg13g2_o21ai_1 _2662_ (.B1(net844),
    .VDD(VPWR),
    .Y(_0870_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_sie.data_q[1] ),
    .A2(_0863_));
 sg13g2_nor2_1 _2663_ (.A(_0864_),
    .B(_0870_),
    .Y(_0871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2664_ (.B1(net601),
    .VDD(VPWR),
    .Y(_0872_),
    .VSS(VGND),
    .A1(net838),
    .A2(_0871_));
 sg13g2_a22oi_1 _2665_ (.Y(_0024_),
    .B1(_0872_),
    .B2(_1973_),
    .A2(_0599_),
    .A1(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2666_ (.Y(_0873_),
    .A(net844),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2667_ (.B1(_0873_),
    .VDD(VPWR),
    .Y(_0025_),
    .VSS(VGND),
    .A1(net141),
    .A2(_0844_));
 sg13g2_nor4_1 _2668_ (.A(net753),
    .B(_0556_),
    .C(_0564_),
    .D(_0585_),
    .Y(_0874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2669_ (.B1(net843),
    .VDD(VPWR),
    .Y(_0875_),
    .VSS(VGND),
    .A1(net598),
    .A2(_0874_));
 sg13g2_o21ai_1 _2670_ (.B1(net1027),
    .VDD(VPWR),
    .Y(_0026_),
    .VSS(VGND),
    .A1(_0572_),
    .A2(_0590_));
 sg13g2_nand2_1 _2671_ (.Y(_0876_),
    .A(net841),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2672_ (.A(net841),
    .B(net524),
    .Y(_0877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2673_ (.B1(_0876_),
    .VDD(VPWR),
    .Y(_0027_),
    .VSS(VGND),
    .A1(_0844_),
    .A2(_0877_));
 sg13g2_nand2_1 _2674_ (.Y(_0878_),
    .A(net838),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2675_ (.B1(_0878_),
    .VDD(VPWR),
    .Y(_0028_),
    .VSS(VGND),
    .A1(_1974_),
    .A2(_0844_));
 sg13g2_a22oi_1 _2676_ (.Y(_0879_),
    .B1(net593),
    .B2(net846),
    .A2(net599),
    .A1(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2677_ (.VDD(VPWR),
    .Y(_0018_),
    .A(net1036),
    .VSS(VGND));
 sg13g2_nand4_1 _2678_ (.B(net710),
    .C(_0511_),
    .A(net841),
    .Y(_0880_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0522_));
 sg13g2_o21ai_1 _2679_ (.B1(_0880_),
    .VDD(VPWR),
    .Y(_0019_),
    .VSS(VGND),
    .A1(_1920_),
    .A2(net601));
 sg13g2_nand2_1 _2680_ (.Y(_0881_),
    .A(net1007),
    .B(_2042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2681_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .Y(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2682_ (.A(_2036_),
    .B(_0882_),
    .Y(_0883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2683_ (.B(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .C(net57),
    .Y(_0884_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ));
 sg13g2_o21ai_1 _2684_ (.B1(_0883_),
    .VDD(VPWR),
    .Y(_0885_),
    .VSS(VGND),
    .A1(_2035_),
    .A2(_0884_));
 sg13g2_nor4_1 _2685_ (.A(_0056_),
    .B(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .C(net312),
    .D(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .Y(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2686_ (.X(_0887_),
    .A(_2036_),
    .B(_2046_),
    .C(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2687_ (.B(_1952_),
    .C(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ),
    .A(_1949_),
    .Y(_0888_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0887_));
 sg13g2_nand3_1 _2688_ (.B(_2036_),
    .C(_0884_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .Y(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2689_ (.B(_0888_),
    .C(_0889_),
    .A(_0885_),
    .Y(_0890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2690_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2038_),
    .A2(_0890_),
    .Y(_0891_),
    .B1(_0881_));
 sg13g2_o21ai_1 _2691_ (.B1(net314),
    .VDD(VPWR),
    .Y(_0892_),
    .VSS(VGND),
    .A1(_1943_),
    .A2(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ));
 sg13g2_a21oi_1 _2692_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net572),
    .A2(net707),
    .Y(_0893_),
    .B1(_0891_));
 sg13g2_o21ai_1 _2693_ (.B1(net573),
    .VDD(VPWR),
    .Y(_0029_),
    .VSS(VGND),
    .A1(_2043_),
    .A2(_0892_));
 sg13g2_nand2b_1 _2694_ (.Y(_0894_),
    .B(_0673_),
    .A_N(_0771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2695_ (.B1(_0894_),
    .VDD(VPWR),
    .Y(_0895_),
    .VSS(VGND),
    .A1(_0650_),
    .A2(_0745_));
 sg13g2_o21ai_1 _2696_ (.B1(net894),
    .VDD(VPWR),
    .Y(_0896_),
    .VSS(VGND),
    .A1(_0812_),
    .A2(_0895_));
 sg13g2_nand3_1 _2697_ (.B(net623),
    .C(_0706_),
    .A(net794),
    .Y(_0897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2698_ (.B1(_0896_),
    .VDD(VPWR),
    .Y(_0002_),
    .VSS(VGND),
    .A1(_0720_),
    .A2(_0897_));
 sg13g2_nand3_1 _2699_ (.B(_2037_),
    .C(_0884_),
    .A(_2032_),
    .Y(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2700_ (.B(_2032_),
    .C(_2037_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .Y(_0899_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0898_));
 sg13g2_inv_1 _2701_ (.VDD(VPWR),
    .Y(_0900_),
    .A(_0899_),
    .VSS(VGND));
 sg13g2_a21oi_2 _2702_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net707),
    .Y(_0901_),
    .A2(_0900_),
    .A1(net976));
 sg13g2_nand2b_1 _2703_ (.Y(_0902_),
    .B(net1007),
    .A_N(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2704_ (.B(_2038_),
    .C(_0884_),
    .A(net1007),
    .Y(_0903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2705_ (.VDD(VPWR),
    .Y(_0904_),
    .A(_0903_),
    .VSS(VGND));
 sg13g2_nand3_1 _2706_ (.B(_0883_),
    .C(_0904_),
    .A(_2042_),
    .Y(_0905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2707_ (.B(net976),
    .C(_2038_),
    .A(net1007),
    .Y(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2708_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2037_),
    .A2(_0882_),
    .Y(_0907_),
    .B1(_0906_));
 sg13g2_nand3_1 _2709_ (.B(_0884_),
    .C(_0907_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .Y(_0908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2710_ (.Y(_0909_),
    .B(_2042_),
    .A_N(_2035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2711_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0910_),
    .B(_2047_),
    .A(_1975_));
 sg13g2_or2_1 _2712_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0911_),
    .B(_0910_),
    .A(_0909_));
 sg13g2_nand4_1 _2713_ (.B(_0905_),
    .C(_0908_),
    .A(_0902_),
    .Y(_0030_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0911_));
 sg13g2_or2_1 _2714_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0912_),
    .B(_2044_),
    .A(_2039_));
 sg13g2_nor3_1 _2715_ (.A(net990),
    .B(_2043_),
    .C(_0429_),
    .Y(_0913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net961),
    .A2(net707),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_nand2_1 _2717_ (.Y(_0031_),
    .A(_0912_),
    .B(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2718_ (.Y(_0915_),
    .A(net314),
    .B(net707),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2719_ (.B1(_0915_),
    .VDD(VPWR),
    .Y(_0032_),
    .VSS(VGND),
    .A1(_0881_),
    .A2(_0888_));
 sg13g2_nor2_1 _2720_ (.A(net717),
    .B(_1976_),
    .Y(_0916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2721_ (.Y(_0917_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .B(_0916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2722_ (.B(net391),
    .C(net457),
    .A(net744),
    .Y(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2723_ (.Y(_0919_),
    .A(net393),
    .B(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2724_ (.B1(net394),
    .VDD(VPWR),
    .Y(_0033_),
    .VSS(VGND),
    .A1(_1977_),
    .A2(_0917_));
 sg13g2_a22oi_1 _2725_ (.Y(_0920_),
    .B1(_0917_),
    .B2(net568),
    .A2(_2006_),
    .A1(net744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2726_ (.VDD(VPWR),
    .Y(_0034_),
    .A(net569),
    .VSS(VGND));
 sg13g2_nor2_1 _2727_ (.A(net393),
    .B(net929),
    .Y(_0921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2728_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1978_),
    .A2(_0918_),
    .Y(_0035_),
    .B1(_0921_));
 sg13g2_nand2_1 _2729_ (.Y(_0922_),
    .A(net308),
    .B(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2730_ (.Y(_0923_),
    .A(net625),
    .B(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2731_ (.A(net626),
    .B(_0923_),
    .Y(_0924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2732_ (.A(net872),
    .B(net924),
    .Y(_0925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2733_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0926_),
    .B(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ));
 sg13g2_a221oi_1 _2734_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1979_),
    .C1(_0925_),
    .B1(_0923_),
    .A1(net625),
    .Y(_0036_),
    .A2(_2028_));
 sg13g2_nand2_1 _2735_ (.Y(_0927_),
    .A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .B(_0923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2736_ (.B1(_0927_),
    .VDD(VPWR),
    .Y(_0037_),
    .VSS(VGND),
    .A1(net368),
    .A2(_2025_));
 sg13g2_a22oi_1 _2737_ (.Y(_0928_),
    .B1(_0924_),
    .B2(net924),
    .A2(_0923_),
    .A1(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2738_ (.VDD(VPWR),
    .Y(_0038_),
    .A(net925),
    .VSS(VGND));
 sg13g2_nand2_1 _2739_ (.Y(_0929_),
    .A(net866),
    .B(_0807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2740_ (.Y(_0930_),
    .A(_0694_),
    .B(_0744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2741_ (.B1(_0929_),
    .VDD(VPWR),
    .Y(_0003_),
    .VSS(VGND),
    .A1(_0632_),
    .A2(_0930_));
 sg13g2_and2_1 _2742_ (.A(net61),
    .B(net49),
    .X(_0041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2743_ (.Y(_0931_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2744_ (.Y(_0932_),
    .A(net813),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2745_ (.Y(_0933_),
    .A(net820),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2746_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .A(net814),
    .X(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2747_ (.B(_0932_),
    .C(_0933_),
    .A(_0931_),
    .Y(_0935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2748_ (.B1(net739),
    .VDD(VPWR),
    .Y(_0936_),
    .VSS(VGND),
    .A1(_0934_),
    .A2(_0935_));
 sg13g2_nand2b_1 _2749_ (.Y(_0937_),
    .B(net543),
    .A_N(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2750_ (.Y(_0042_),
    .A(_0936_),
    .B(_0937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2751_ (.Y(_0938_),
    .A(net532),
    .B(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2752_ (.Y(_0939_),
    .A(net452),
    .B(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2753_ (.Y(_0940_),
    .A(_0938_),
    .B(_0939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2754_ (.A(net53),
    .B(_0940_),
    .Y(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2755_ (.Y(_0941_),
    .B(net567),
    .A_N(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2756_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net708),
    .A2(_0941_),
    .Y(_0047_),
    .B1(_0940_));
 sg13g2_or2_1 _2757_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0942_),
    .B(_0908_),
    .A(net707));
 sg13g2_nor2b_1 _2758_ (.A(net450),
    .B_N(net614),
    .Y(_0943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2759_ (.A(net748),
    .B(_0943_),
    .Y(_0045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2760_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ),
    .A2(_2042_),
    .Y(_0944_),
    .B1(net305));
 sg13g2_nor2_1 _2761_ (.A(net748),
    .B(net306),
    .Y(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2762_ (.A(net501),
    .B_N(_2049_),
    .Y(_0945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2763_ (.A(net748),
    .B(net502),
    .Y(_0043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2764_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1909_),
    .Y(net28),
    .A2(_1993_),
    .A1(net835));
 sg13g2_a21oi_1 _2765_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .A2(_1993_),
    .Y(net30),
    .B1(_0054_));
 sg13g2_xor2_1 _2766_ (.B(net49),
    .A(net61),
    .X(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2767_ (.A(\u_usb_cdc.bus_reset ),
    .B_N(net726),
    .Y(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2768_ (.Y(_0946_),
    .B(_0452_),
    .A_N(_0450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2769_ (.A2(_0946_),
    .A1(_0479_),
    .B1(_0441_),
    .X(_0947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2770_ (.B(_0450_),
    .C(_0479_),
    .A(net838),
    .Y(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2771_ (.X(_0949_),
    .A(_0841_),
    .B(_0947_),
    .C(_0948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2772_ (.A(net840),
    .B(net839),
    .Y(_0950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2773_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0951_),
    .B(net839),
    .A(net840));
 sg13g2_nand4_1 _2774_ (.B(_0522_),
    .C(_0949_),
    .A(_0512_),
    .Y(_0952_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0951_));
 sg13g2_nand2_1 _2775_ (.Y(_0953_),
    .A(net769),
    .B(\u_usb_cdc.u_sie.out_toggle_q[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2776_ (.B1(_0953_),
    .VDD(VPWR),
    .Y(_0954_),
    .VSS(VGND),
    .A1(net769),
    .A2(_1987_));
 sg13g2_xnor2_1 _2777_ (.Y(_0955_),
    .A(\u_usb_cdc.u_sie.pid_q[3] ),
    .B(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2778_ (.Y(_0956_),
    .A(net710),
    .B(_0955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2779_ (.A(net768),
    .B(_0952_),
    .C(_0956_),
    .Y(_0957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2780_ (.A(net486),
    .B(_0957_),
    .Y(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2781_ (.A(net840),
    .B(_0952_),
    .Y(_0959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2782_ (.A(net768),
    .B(_1987_),
    .C(_0952_),
    .D(_0956_),
    .Y(_0960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2783_ (.A(_0958_),
    .B(_0959_),
    .C(_0960_),
    .Y(_0067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2784_ (.A(net850),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .C(_0551_),
    .D(_0747_),
    .Y(_0961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2785_ (.A(\u_usb_cdc.u_ctrl_endp.endp_q[1] ),
    .B(_1970_),
    .C(net545),
    .D(net500),
    .Y(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2786_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1971_),
    .A2(_0962_),
    .Y(_0963_),
    .B1(net851));
 sg13g2_nor2b_2 _2787_ (.A(_0963_),
    .B_N(_0961_),
    .Y(_0964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2788_ (.Y(_0965_),
    .A(net742),
    .B(_0964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2789_ (.B(net638),
    .C(_0955_),
    .Y(_0966_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net771));
 sg13g2_nor2_1 _2790_ (.A(net752),
    .B(_0964_),
    .Y(_0967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2791_ (.Y(_0968_),
    .A(_0438_),
    .B(_0967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2792_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net840),
    .A2(_0513_),
    .Y(_0969_),
    .B1(_0968_));
 sg13g2_a22oi_1 _2793_ (.Y(_0970_),
    .B1(_0964_),
    .B2(net745),
    .A2(_0600_),
    .A1(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2794_ (.A(_0966_),
    .B(_0969_),
    .C(_0970_),
    .Y(_0971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2795_ (.B1(_0965_),
    .VDD(VPWR),
    .Y(_0972_),
    .VSS(VGND),
    .A1(net55),
    .A2(_0971_));
 sg13g2_a21oi_1 _2796_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net55),
    .A2(_0971_),
    .Y(_0068_),
    .B1(_0972_));
 sg13g2_nand2_1 _2797_ (.Y(_0973_),
    .A(net560),
    .B(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2798_ (.A(net767),
    .B(_0973_),
    .Y(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2799_ (.B1(net750),
    .VDD(VPWR),
    .Y(_0975_),
    .VSS(VGND),
    .A1(net839),
    .A2(_0974_));
 sg13g2_o21ai_1 _2800_ (.B1(_0975_),
    .VDD(VPWR),
    .Y(_0976_),
    .VSS(VGND),
    .A1(net839),
    .A2(net844));
 sg13g2_nor4_1 _2801_ (.A(net519),
    .B(\u_usb_cdc.u_sie.data_q[3] ),
    .C(_2017_),
    .D(_0854_),
    .Y(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2802_ (.Y(_0978_),
    .A(_0974_),
    .B(_0977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2803_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net844),
    .A2(_0978_),
    .Y(_0979_),
    .B1(_0976_));
 sg13g2_nand3_1 _2804_ (.B(_0949_),
    .C(_0979_),
    .A(net593),
    .Y(_0980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2805_ (.B1(net406),
    .VDD(VPWR),
    .Y(_0981_),
    .VSS(VGND),
    .A1(_0516_),
    .A2(_0980_));
 sg13g2_nand2_1 _2806_ (.Y(_0982_),
    .A(\u_usb_cdc.u_sie.in_toggle_q[1] ),
    .B(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2807_ (.A(net768),
    .B_N(\u_usb_cdc.endp[1] ),
    .Y(_0983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2808_ (.Y(_0984_),
    .B1(_0983_),
    .B2(\u_usb_cdc.u_sie.in_toggle_q[2] ),
    .A2(_0514_),
    .A1(\u_usb_cdc.u_sie.in_toggle_q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2809_ (.A(net768),
    .B(\u_usb_cdc.endp[1] ),
    .C(net406),
    .D(_2014_),
    .Y(_0985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2810_ (.A(net838),
    .B(_0985_),
    .Y(_0986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2811_ (.B1(_0981_),
    .VDD(VPWR),
    .Y(_0069_),
    .VSS(VGND),
    .A1(_0980_),
    .A2(_0986_));
 sg13g2_nor2_1 _2812_ (.A(_0523_),
    .B(_0978_),
    .Y(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2813_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0988_),
    .B(_0978_),
    .A(_0523_));
 sg13g2_nand2_1 _2814_ (.Y(_0989_),
    .A(net638),
    .B(_0987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2815_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2014_),
    .Y(_0990_),
    .A2(_0984_),
    .A1(_0982_));
 sg13g2_nor2b_1 _2816_ (.A(_0514_),
    .B_N(\u_usb_cdc.endp[3] ),
    .Y(_0991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2817_ (.A(\u_usb_cdc.endp[2] ),
    .B(_0988_),
    .C(_0990_),
    .D(_0991_),
    .Y(_0992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2818_ (.Y(_0993_),
    .B1(_0992_),
    .B2(_0566_),
    .A2(_0989_),
    .A1(net856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _2819_ (.A2(_0962_),
    .A1(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .B1(net851),
    .X(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2820_ (.A(net742),
    .B(_0961_),
    .X(_0995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2821_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0994_),
    .A2(_0995_),
    .Y(_0070_),
    .B1(net857));
 sg13g2_nor2b_1 _2822_ (.A(_2014_),
    .B_N(_0983_),
    .Y(_0996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2823_ (.Y(_0997_),
    .A(_0987_),
    .B(_0996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2824_ (.Y(_0998_),
    .B1(_0997_),
    .B2(net378),
    .A2(_0992_),
    .A1(_0983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2825_ (.Y(_0999_),
    .A(\u_usb_cdc.u_ctrl_endp.endp_q[1] ),
    .B(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _2826_ (.A(\u_usb_cdc.u_ctrl_endp.endp_q[0] ),
    .B(\u_usb_cdc.u_ctrl_endp.endp_q[2] ),
    .C(\u_usb_cdc.u_ctrl_endp.endp_q[3] ),
    .D(_0999_),
    .Y(_1000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2827_ (.B1(_0995_),
    .VDD(VPWR),
    .Y(_1001_),
    .VSS(VGND),
    .A1(net851),
    .A2(_1000_));
 sg13g2_nor2b_1 _2828_ (.A(net379),
    .B_N(_1001_),
    .Y(_0071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _2829_ (.X(_1002_),
    .A(net838),
    .B(_0479_),
    .C(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2830_ (.B(\u_usb_cdc.addr[0] ),
    .C(net594),
    .A(net838),
    .Y(_1003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2831_ (.Y(_1004_),
    .B(_1003_),
    .A_N(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _2832_ (.B(_0479_),
    .C(net763),
    .Y(_1005_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net750));
 sg13g2_a21oi_1 _2833_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net838),
    .A2(net594),
    .Y(_1006_),
    .B1(net261));
 sg13g2_a21oi_1 _2834_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1004_),
    .A2(_1005_),
    .Y(_0072_),
    .B1(net262));
 sg13g2_nand2_1 _2835_ (.Y(_1007_),
    .A(net299),
    .B(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _2836_ (.A(net835),
    .B(_0926_),
    .Y(_1008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _2837_ (.A(net626),
    .B_N(_1008_),
    .Y(_1009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2838_ (.Y(_1010_),
    .B(_1008_),
    .A_N(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2839_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .C1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .B1(_2028_),
    .A1(_1909_),
    .Y(_1011_),
    .A2(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ));
 sg13g2_a21oi_1 _2840_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1010_),
    .A2(_1011_),
    .Y(_1012_),
    .B1(_2022_));
 sg13g2_a22oi_1 _2841_ (.Y(_1013_),
    .B1(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .B2(net625),
    .A2(net747),
    .A1(_1909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2842_ (.B1(_1007_),
    .VDD(VPWR),
    .Y(_0073_),
    .VSS(VGND),
    .A1(_1012_),
    .A2(_1013_));
 sg13g2_nand2_1 _2843_ (.Y(_1014_),
    .A(net933),
    .B(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2844_ (.Y(_1015_),
    .A(net834),
    .B(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2845_ (.B(net833),
    .C(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .A(net977),
    .Y(_1016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2846_ (.A(_1985_),
    .B(_1016_),
    .Y(_1017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2847_ (.A(net834),
    .B(net833),
    .Y(_1018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _2848_ (.A(net834),
    .B(net833),
    .C(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .Y(_1019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2849_ (.Y(_1020_),
    .B(net994),
    .A_N(_1019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1016_),
    .A2(_1020_),
    .Y(_1021_),
    .B1(_1017_));
 sg13g2_xor2_1 _2851_ (.B(_1021_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .X(_1022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _2852_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net834),
    .Y(_1023_),
    .A2(_1019_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ));
 sg13g2_xnor2_1 _2853_ (.Y(_1024_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .B(_1023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2854_ (.B(net1044),
    .A(net977),
    .X(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2855_ (.Y(_1026_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .A_N(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2856_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1986_),
    .A2(_1025_),
    .Y(_1027_),
    .B1(_1017_));
 sg13g2_xnor2_1 _2857_ (.Y(_1028_),
    .A(net1025),
    .B(_1015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _2858_ (.Y(_1029_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .B(_1028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _2859_ (.B(_1026_),
    .C(_1027_),
    .A(_1024_),
    .Y(_1030_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1029_));
 sg13g2_o21ai_1 _2860_ (.B1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ),
    .VDD(VPWR),
    .Y(_1031_),
    .VSS(VGND),
    .A1(_1022_),
    .A2(_1030_));
 sg13g2_or2_1 _2861_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1032_),
    .B(_1031_),
    .A(net716));
 sg13g2_nand2_2 _2862_ (.Y(_1033_),
    .A(net547),
    .B(_1032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2863_ (.Y(_0074_),
    .A(net647),
    .B(_1033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2864_ (.A0(net2),
    .A1(net1018),
    .S(net646),
    .X(_0075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2865_ (.A0(net3),
    .A1(net1013),
    .S(net646),
    .X(_0076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2866_ (.A0(net4),
    .A1(net1006),
    .S(net646),
    .X(_0077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2867_ (.A0(net5),
    .A1(net996),
    .S(net646),
    .X(_0078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2868_ (.A0(net6),
    .A1(net1000),
    .S(net646),
    .X(_0079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2869_ (.A0(net7),
    .A1(net1002),
    .S(net646),
    .X(_0080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2870_ (.A0(net8),
    .A1(net1010),
    .S(net646),
    .X(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2871_ (.A0(net9),
    .A1(net1020),
    .S(net646),
    .X(_0082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _2872_ (.A(net833),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .C(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .Y(_1034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2873_ (.A(_1985_),
    .B(_1019_),
    .X(_1035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2874_ (.Y(_1036_),
    .A(net740),
    .B(_1035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2875_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .A1(net461),
    .S(_1036_),
    .X(_0083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2876_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .A1(net549),
    .S(_1036_),
    .X(_0084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2877_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .A1(net490),
    .S(_1036_),
    .X(_0085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2878_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .A1(net433),
    .S(_1036_),
    .X(_0086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2879_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .A1(net443),
    .S(_1036_),
    .X(_0087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2880_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .A1(net455),
    .S(_1036_),
    .X(_0088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2881_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .A1(net526),
    .S(_1036_),
    .X(_0089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2882_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .A1(net869),
    .S(_1036_),
    .X(_0090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2883_ (.B(net834),
    .C(_1034_),
    .A(net740),
    .Y(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2884_ (.Y(_1038_),
    .A(net82),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2885_ (.A(net833),
    .B_N(net834),
    .Y(_1039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2886_ (.Y(_1040_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _2887_ (.B(_1018_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .X(_1041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2888_ (.Y(_1042_),
    .A(net740),
    .B(_1020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2889_ (.A(_1035_),
    .B(_1042_),
    .Y(_1043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2890_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1044_),
    .B(_1042_),
    .A(_1041_));
 sg13g2_o21ai_1 _2891_ (.B1(_1038_),
    .VDD(VPWR),
    .Y(_0091_),
    .VSS(VGND),
    .A1(_1040_),
    .A2(net620));
 sg13g2_nand2_1 _2892_ (.Y(_1045_),
    .A(net193),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2893_ (.Y(_1046_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2894_ (.B1(_1045_),
    .VDD(VPWR),
    .Y(_0092_),
    .VSS(VGND),
    .A1(net618),
    .A2(_1046_));
 sg13g2_nand2_1 _2895_ (.Y(_1047_),
    .A(net76),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2896_ (.Y(_1048_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2897_ (.B1(_1047_),
    .VDD(VPWR),
    .Y(_0093_),
    .VSS(VGND),
    .A1(net618),
    .A2(_1048_));
 sg13g2_nand2_1 _2898_ (.Y(_1049_),
    .A(net78),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2899_ (.Y(_1050_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2900_ (.B1(_1049_),
    .VDD(VPWR),
    .Y(_0094_),
    .VSS(VGND),
    .A1(net618),
    .A2(_1050_));
 sg13g2_nand2_1 _2901_ (.Y(_1051_),
    .A(net119),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2902_ (.Y(_1052_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2903_ (.B1(_1051_),
    .VDD(VPWR),
    .Y(_0095_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1052_));
 sg13g2_nand2_1 _2904_ (.Y(_1053_),
    .A(net131),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2905_ (.Y(_1054_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2906_ (.B1(_1053_),
    .VDD(VPWR),
    .Y(_0096_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1054_));
 sg13g2_nand2_1 _2907_ (.Y(_1055_),
    .A(net220),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2908_ (.Y(_1056_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .B(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2909_ (.B1(_1055_),
    .VDD(VPWR),
    .Y(_0097_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1056_));
 sg13g2_nand2_1 _2910_ (.Y(_1057_),
    .A(net105),
    .B(_1037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2911_ (.Y(_1058_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .B(_1039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2912_ (.B1(_1057_),
    .VDD(VPWR),
    .Y(_0098_),
    .VSS(VGND),
    .A1(net620),
    .A2(_1058_));
 sg13g2_nor2b_2 _2913_ (.A(net834),
    .B_N(net833),
    .Y(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2914_ (.Y(_1060_),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net618));
 sg13g2_nand2_1 _2915_ (.Y(_1061_),
    .A(net250),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2916_ (.Y(_1062_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2917_ (.B1(_1061_),
    .VDD(VPWR),
    .Y(_0099_),
    .VSS(VGND),
    .A1(net620),
    .A2(_1062_));
 sg13g2_nand2_1 _2918_ (.Y(_1063_),
    .A(net168),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2919_ (.Y(_1064_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2920_ (.B1(_1063_),
    .VDD(VPWR),
    .Y(_0100_),
    .VSS(VGND),
    .A1(net618),
    .A2(_1064_));
 sg13g2_nand2_1 _2921_ (.Y(_1065_),
    .A(net182),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2922_ (.Y(_1066_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2923_ (.B1(_1065_),
    .VDD(VPWR),
    .Y(_0101_),
    .VSS(VGND),
    .A1(net618),
    .A2(_1066_));
 sg13g2_nand2_1 _2924_ (.Y(_1067_),
    .A(net248),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2925_ (.Y(_1068_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2926_ (.B1(_1067_),
    .VDD(VPWR),
    .Y(_0102_),
    .VSS(VGND),
    .A1(net618),
    .A2(_1068_));
 sg13g2_nand2_1 _2927_ (.Y(_1069_),
    .A(net94),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2928_ (.Y(_1070_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2929_ (.B1(_1069_),
    .VDD(VPWR),
    .Y(_0103_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1070_));
 sg13g2_nand2_1 _2930_ (.Y(_1071_),
    .A(net72),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2931_ (.Y(_1072_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .B(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2932_ (.B1(_1071_),
    .VDD(VPWR),
    .Y(_0104_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1072_));
 sg13g2_nand2_1 _2933_ (.Y(_1073_),
    .A(net238),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2934_ (.Y(_1074_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .B(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2935_ (.B1(_1073_),
    .VDD(VPWR),
    .Y(_0105_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1074_));
 sg13g2_nand2_1 _2936_ (.Y(_1075_),
    .A(net121),
    .B(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2937_ (.Y(_1076_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .B(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2938_ (.B1(_1075_),
    .VDD(VPWR),
    .Y(_0106_),
    .VSS(VGND),
    .A1(net621),
    .A2(_1076_));
 sg13g2_nor2_2 _2939_ (.A(_1015_),
    .B(net621),
    .Y(_1077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2940_ (.A0(net515),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .S(_1077_),
    .X(_0107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2941_ (.A0(net511),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .S(_1077_),
    .X(_0108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2942_ (.A0(net537),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .S(_1077_),
    .X(_0109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2943_ (.A0(net528),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .S(_1077_),
    .X(_0110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2944_ (.A0(net535),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .S(_1077_),
    .X(_0111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2945_ (.A0(net520),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .S(_1077_),
    .X(_0112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2946_ (.A0(net570),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .S(_1077_),
    .X(_0113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _2947_ (.A0(net509),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .S(_1077_),
    .X(_0114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2948_ (.A(_1034_),
    .B_N(_1018_),
    .Y(_1078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _2949_ (.Y(_1079_),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net620));
 sg13g2_nand2_1 _2950_ (.Y(_1080_),
    .A(net158),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2951_ (.Y(_1081_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .B(_1078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2952_ (.B1(_1080_),
    .VDD(VPWR),
    .Y(_0115_),
    .VSS(VGND),
    .A1(net620),
    .A2(_1081_));
 sg13g2_nand2_1 _2953_ (.Y(_1082_),
    .A(net218),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2954_ (.Y(_1083_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2955_ (.B1(_1082_),
    .VDD(VPWR),
    .Y(_0116_),
    .VSS(VGND),
    .A1(net620),
    .A2(_1083_));
 sg13g2_nand2_1 _2956_ (.Y(_1084_),
    .A(net154),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2957_ (.Y(_1085_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2958_ (.B1(_1084_),
    .VDD(VPWR),
    .Y(_0117_),
    .VSS(VGND),
    .A1(net620),
    .A2(_1085_));
 sg13g2_nand2_1 _2959_ (.Y(_1086_),
    .A(net198),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2960_ (.Y(_1087_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2961_ (.B1(_1086_),
    .VDD(VPWR),
    .Y(_0118_),
    .VSS(VGND),
    .A1(net618),
    .A2(_1087_));
 sg13g2_nand2_1 _2962_ (.Y(_1088_),
    .A(net205),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2963_ (.Y(_1089_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2964_ (.B1(_1088_),
    .VDD(VPWR),
    .Y(_0119_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1089_));
 sg13g2_nand2_1 _2965_ (.Y(_1090_),
    .A(net113),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2966_ (.Y(_1091_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2967_ (.B1(_1090_),
    .VDD(VPWR),
    .Y(_0120_),
    .VSS(VGND),
    .A1(net619),
    .A2(_1091_));
 sg13g2_nand2_1 _2968_ (.Y(_1092_),
    .A(net196),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2969_ (.Y(_1093_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2970_ (.B1(_1092_),
    .VDD(VPWR),
    .Y(_0121_),
    .VSS(VGND),
    .A1(net621),
    .A2(_1093_));
 sg13g2_nand2_1 _2971_ (.Y(_1094_),
    .A(net177),
    .B(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2972_ (.Y(_1095_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .B(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2973_ (.B1(_1094_),
    .VDD(VPWR),
    .Y(_0122_),
    .VSS(VGND),
    .A1(net620),
    .A2(_1095_));
 sg13g2_nand4_1 _2974_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .C(_1985_),
    .A(net740),
    .Y(_1096_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net645));
 sg13g2_nand2_1 _2975_ (.Y(_1097_),
    .A(net62),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _2976_ (.Y(_1098_),
    .A(net740),
    .B(_1041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2977_ (.Y(_1099_),
    .A(_1041_),
    .B(_1043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2978_ (.VDD(VPWR),
    .Y(_1100_),
    .A(net610),
    .VSS(VGND));
 sg13g2_o21ai_1 _2979_ (.B1(_1097_),
    .VDD(VPWR),
    .Y(_0123_),
    .VSS(VGND),
    .A1(_1040_),
    .A2(net612));
 sg13g2_nand2_1 _2980_ (.Y(_1101_),
    .A(net64),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2981_ (.B1(_1101_),
    .VDD(VPWR),
    .Y(_0124_),
    .VSS(VGND),
    .A1(_1046_),
    .A2(net610));
 sg13g2_nand2_1 _2982_ (.Y(_1102_),
    .A(net74),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2983_ (.B1(_1102_),
    .VDD(VPWR),
    .Y(_0125_),
    .VSS(VGND),
    .A1(_1048_),
    .A2(net610));
 sg13g2_nand2_1 _2984_ (.Y(_1103_),
    .A(net59),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2985_ (.B1(_1103_),
    .VDD(VPWR),
    .Y(_0126_),
    .VSS(VGND),
    .A1(_1050_),
    .A2(net610));
 sg13g2_nand2_1 _2986_ (.Y(_1104_),
    .A(net90),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2987_ (.B1(_1104_),
    .VDD(VPWR),
    .Y(_0127_),
    .VSS(VGND),
    .A1(_1052_),
    .A2(net610));
 sg13g2_nand2_1 _2988_ (.Y(_1105_),
    .A(net117),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2989_ (.B1(_1105_),
    .VDD(VPWR),
    .Y(_0128_),
    .VSS(VGND),
    .A1(_1054_),
    .A2(net611));
 sg13g2_nand2_1 _2990_ (.Y(_1106_),
    .A(net70),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2991_ (.B1(_1106_),
    .VDD(VPWR),
    .Y(_0129_),
    .VSS(VGND),
    .A1(_1056_),
    .A2(net611));
 sg13g2_nand2_1 _2992_ (.Y(_1107_),
    .A(net96),
    .B(_1096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2993_ (.B1(_1107_),
    .VDD(VPWR),
    .Y(_0130_),
    .VSS(VGND),
    .A1(_1058_),
    .A2(net612));
 sg13g2_nand2_2 _2994_ (.Y(_1108_),
    .A(net644),
    .B(_1100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2995_ (.Y(_1109_),
    .A(net88),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2996_ (.B1(_1109_),
    .VDD(VPWR),
    .Y(_0131_),
    .VSS(VGND),
    .A1(_1062_),
    .A2(net612));
 sg13g2_nand2_1 _2997_ (.Y(_1110_),
    .A(net80),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2998_ (.B1(_1110_),
    .VDD(VPWR),
    .Y(_0132_),
    .VSS(VGND),
    .A1(_1064_),
    .A2(net610));
 sg13g2_nand2_1 _2999_ (.Y(_1111_),
    .A(net253),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3000_ (.B1(_1111_),
    .VDD(VPWR),
    .Y(_0133_),
    .VSS(VGND),
    .A1(_1066_),
    .A2(net610));
 sg13g2_nand2_1 _3001_ (.Y(_1112_),
    .A(net86),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3002_ (.B1(_1112_),
    .VDD(VPWR),
    .Y(_0134_),
    .VSS(VGND),
    .A1(_1068_),
    .A2(net610));
 sg13g2_nand2_1 _3003_ (.Y(_1113_),
    .A(net135),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3004_ (.B1(_1113_),
    .VDD(VPWR),
    .Y(_0135_),
    .VSS(VGND),
    .A1(_1070_),
    .A2(net611));
 sg13g2_nand2_1 _3005_ (.Y(_1114_),
    .A(net240),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3006_ (.B1(_1114_),
    .VDD(VPWR),
    .Y(_0136_),
    .VSS(VGND),
    .A1(_1072_),
    .A2(net611));
 sg13g2_nand2_1 _3007_ (.Y(_1115_),
    .A(net242),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3008_ (.B1(_1115_),
    .VDD(VPWR),
    .Y(_0137_),
    .VSS(VGND),
    .A1(_1074_),
    .A2(net611));
 sg13g2_nand2_1 _3009_ (.Y(_1116_),
    .A(net150),
    .B(_1108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3010_ (.B1(_1116_),
    .VDD(VPWR),
    .Y(_0138_),
    .VSS(VGND),
    .A1(_1076_),
    .A2(net612));
 sg13g2_or2_1 _3011_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1117_),
    .B(net612),
    .A(_1015_));
 sg13g2_mux2_1 _3012_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .A1(net507),
    .S(_1117_),
    .X(_0139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3013_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .A1(net517),
    .S(_1117_),
    .X(_0140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3014_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .A1(net469),
    .S(_1117_),
    .X(_0141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3015_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .A1(net467),
    .S(_1117_),
    .X(_0142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3016_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .A1(net475),
    .S(_1117_),
    .X(_0143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3017_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .A1(net463),
    .S(_1117_),
    .X(_0144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3018_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .A1(net479),
    .S(_1117_),
    .X(_0145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3019_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .A1(net477),
    .S(_1117_),
    .X(_0146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3020_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .C(_1019_),
    .A(net740),
    .Y(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3021_ (.Y(_1119_),
    .A(net92),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3022_ (.B1(_1119_),
    .VDD(VPWR),
    .Y(_0147_),
    .VSS(VGND),
    .A1(_1081_),
    .A2(_1098_));
 sg13g2_nand2_1 _3023_ (.Y(_1120_),
    .A(net200),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3024_ (.B1(_1120_),
    .VDD(VPWR),
    .Y(_0148_),
    .VSS(VGND),
    .A1(_1083_),
    .A2(_1098_));
 sg13g2_nand2_1 _3025_ (.Y(_1121_),
    .A(net109),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3026_ (.B1(_1121_),
    .VDD(VPWR),
    .Y(_0149_),
    .VSS(VGND),
    .A1(_1085_),
    .A2(_1098_));
 sg13g2_nand2_1 _3027_ (.Y(_1122_),
    .A(net123),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3028_ (.B1(_1122_),
    .VDD(VPWR),
    .Y(_0150_),
    .VSS(VGND),
    .A1(_1087_),
    .A2(_1098_));
 sg13g2_nand2_1 _3029_ (.Y(_1123_),
    .A(net133),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3030_ (.B1(_1123_),
    .VDD(VPWR),
    .Y(_0151_),
    .VSS(VGND),
    .A1(_1089_),
    .A2(_1098_));
 sg13g2_nand2_1 _3031_ (.Y(_1124_),
    .A(net139),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3032_ (.B1(_1124_),
    .VDD(VPWR),
    .Y(_0152_),
    .VSS(VGND),
    .A1(_1091_),
    .A2(_1098_));
 sg13g2_nand2_1 _3033_ (.Y(_1125_),
    .A(net68),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3034_ (.B1(_1125_),
    .VDD(VPWR),
    .Y(_0153_),
    .VSS(VGND),
    .A1(_1093_),
    .A2(_1098_));
 sg13g2_nand2_1 _3035_ (.Y(_1126_),
    .A(net137),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3036_ (.B1(_1126_),
    .VDD(VPWR),
    .Y(_0154_),
    .VSS(VGND),
    .A1(_1095_),
    .A2(_1098_));
 sg13g2_nand2_1 _3037_ (.Y(_1127_),
    .A(net742),
    .B(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3038_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1127_),
    .Y(_1128_),
    .A2(_0593_),
    .A1(_0592_));
 sg13g2_mux2_1 _3039_ (.A0(_1025_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .S(_1031_),
    .X(_1129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3040_ (.A0(net859),
    .A1(_1129_),
    .S(_1128_),
    .X(_0155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3041_ (.A0(_1028_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .S(_1031_),
    .X(_1130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3042_ (.A0(net862),
    .A1(_1130_),
    .S(_1128_),
    .X(_0156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3043_ (.A0(_1021_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .S(_1031_),
    .X(_1131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3044_ (.A0(net882),
    .A1(_1131_),
    .S(_1128_),
    .X(_0157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3045_ (.B1(net647),
    .VDD(VPWR),
    .Y(_1132_),
    .VSS(VGND),
    .A1(net933),
    .A2(_1033_));
 sg13g2_inv_1 _3046_ (.VDD(VPWR),
    .Y(_0158_),
    .A(_1132_),
    .VSS(VGND));
 sg13g2_mux2_1 _3047_ (.A0(_1023_),
    .A1(net977),
    .S(_1032_),
    .X(_0159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3048_ (.A0(_1025_),
    .A1(net833),
    .S(_1032_),
    .X(_0160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3049_ (.A0(_1028_),
    .A1(net1025),
    .S(_1032_),
    .X(_0161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3050_ (.A0(_1021_),
    .A1(net994),
    .S(_1032_),
    .X(_0162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3051_ (.Y(_1133_),
    .A(net1034),
    .B(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3052_ (.Y(_1134_),
    .A(net1037),
    .B(_1133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3053_ (.B(_1128_),
    .C(_1133_),
    .A(\u_usb_cdc.sie_in_data_ack ),
    .Y(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3054_ (.A0(net809),
    .A1(net931),
    .S(_1135_),
    .X(_0163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3055_ (.A(net801),
    .B(_1135_),
    .Y(_1136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3056_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1986_),
    .A2(_1135_),
    .Y(_0164_),
    .B1(_1136_));
 sg13g2_nand2_1 _3057_ (.Y(_1137_),
    .A(net419),
    .B(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3058_ (.B1(_1137_),
    .VDD(VPWR),
    .Y(_0165_),
    .VSS(VGND),
    .A1(_1923_),
    .A2(_1135_));
 sg13g2_nand2_1 _3059_ (.Y(_1138_),
    .A(net363),
    .B(_1135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3060_ (.B1(_1138_),
    .VDD(VPWR),
    .Y(_0166_),
    .VSS(VGND),
    .A1(_1924_),
    .A2(_1135_));
 sg13g2_nor2_1 _3061_ (.A(net829),
    .B(net826),
    .Y(_1139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3062_ (.A(net829),
    .B(net827),
    .C(net826),
    .Y(_1140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3063_ (.Y(_1141_),
    .A(net711),
    .B(_1139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3064_ (.B(_1140_),
    .C(net739),
    .Y(_1142_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net831));
 sg13g2_nand2_1 _3065_ (.Y(_1143_),
    .A(net216),
    .B(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3066_ (.B1(_1143_),
    .VDD(VPWR),
    .Y(_0167_),
    .VSS(VGND),
    .A1(net723),
    .A2(net634));
 sg13g2_nand2_1 _3067_ (.Y(_1144_),
    .A(net252),
    .B(_1142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3068_ (.B1(_1144_),
    .VDD(VPWR),
    .Y(_0168_),
    .VSS(VGND),
    .A1(net722),
    .A2(net635));
 sg13g2_nand2_1 _3069_ (.Y(_1145_),
    .A(net288),
    .B(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3070_ (.B1(_1145_),
    .VDD(VPWR),
    .Y(_0169_),
    .VSS(VGND),
    .A1(_1913_),
    .A2(net634));
 sg13g2_nand2_1 _3071_ (.Y(_1146_),
    .A(net184),
    .B(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3072_ (.B1(_1146_),
    .VDD(VPWR),
    .Y(_0170_),
    .VSS(VGND),
    .A1(net720),
    .A2(net635));
 sg13g2_nand2_1 _3073_ (.Y(_1147_),
    .A(net304),
    .B(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3074_ (.B1(_1147_),
    .VDD(VPWR),
    .Y(_0171_),
    .VSS(VGND),
    .A1(_1915_),
    .A2(net634));
 sg13g2_nand2_1 _3075_ (.Y(_1148_),
    .A(net286),
    .B(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3076_ (.B1(_1148_),
    .VDD(VPWR),
    .Y(_0172_),
    .VSS(VGND),
    .A1(_1914_),
    .A2(net634));
 sg13g2_nand2_1 _3077_ (.Y(_1149_),
    .A(net255),
    .B(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3078_ (.B1(_1149_),
    .VDD(VPWR),
    .Y(_0173_),
    .VSS(VGND),
    .A1(_1917_),
    .A2(net635));
 sg13g2_nand2_1 _3079_ (.Y(_1150_),
    .A(net202),
    .B(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3080_ (.B1(_1150_),
    .VDD(VPWR),
    .Y(_0174_),
    .VSS(VGND),
    .A1(net719),
    .A2(net635));
 sg13g2_nand3_1 _3081_ (.B(net831),
    .C(_1140_),
    .A(net739),
    .Y(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3082_ (.Y(_1152_),
    .A(net203),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3083_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1153_),
    .B(net829),
    .A(net830));
 sg13g2_nor2_2 _3084_ (.A(net827),
    .B(_1153_),
    .Y(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3085_ (.Y(_1155_),
    .A(net739),
    .B(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3086_ (.B(net826),
    .C(_1154_),
    .A(net739),
    .Y(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3087_ (.Y(_1157_),
    .A(net826),
    .B(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3088_ (.Y(_1158_),
    .A(net739),
    .B(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3089_ (.A(net829),
    .B(_1158_),
    .Y(_1159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3090_ (.B(net832),
    .C(_1159_),
    .A(net764),
    .Y(_1160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3091_ (.B1(_1152_),
    .VDD(VPWR),
    .Y(_0175_),
    .VSS(VGND),
    .A1(net828),
    .A2(_1160_));
 sg13g2_nand2_1 _3092_ (.Y(_1161_),
    .A(net103),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3093_ (.B(net832),
    .C(_1159_),
    .A(net762),
    .Y(_1162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3094_ (.B1(_1161_),
    .VDD(VPWR),
    .Y(_0176_),
    .VSS(VGND),
    .A1(net828),
    .A2(_1162_));
 sg13g2_nand2_1 _3095_ (.Y(_1163_),
    .A(net66),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3096_ (.B(net832),
    .C(_1159_),
    .A(net761),
    .Y(_1164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3097_ (.B1(_1163_),
    .VDD(VPWR),
    .Y(_0177_),
    .VSS(VGND),
    .A1(net828),
    .A2(_1164_));
 sg13g2_nand2_1 _3098_ (.Y(_1165_),
    .A(net278),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3099_ (.B(net830),
    .C(_1159_),
    .A(net760),
    .Y(_1166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3100_ (.B1(_1165_),
    .VDD(VPWR),
    .Y(_0178_),
    .VSS(VGND),
    .A1(net827),
    .A2(_1166_));
 sg13g2_nand2_1 _3101_ (.Y(_1167_),
    .A(net111),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3102_ (.B(net832),
    .C(_1159_),
    .A(net759),
    .Y(_1168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3103_ (.B1(_1167_),
    .VDD(VPWR),
    .Y(_0179_),
    .VSS(VGND),
    .A1(net828),
    .A2(_1168_));
 sg13g2_nand2_1 _3104_ (.Y(_1169_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3105_ (.B(net832),
    .C(_1159_),
    .A(\u_usb_cdc.sie_out_data[5] ),
    .Y(_1170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3106_ (.B1(_1169_),
    .VDD(VPWR),
    .Y(_0180_),
    .VSS(VGND),
    .A1(net268),
    .A2(_1170_));
 sg13g2_nand2_1 _3107_ (.Y(_1171_),
    .A(net222),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3108_ (.B(net830),
    .C(_1159_),
    .A(net758),
    .Y(_1172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3109_ (.B1(_1171_),
    .VDD(VPWR),
    .Y(_0181_),
    .VSS(VGND),
    .A1(net827),
    .A2(_1172_));
 sg13g2_nand2_1 _3110_ (.Y(_1173_),
    .A(net115),
    .B(_1151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3111_ (.B(net832),
    .C(_1159_),
    .A(net757),
    .Y(_1174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3112_ (.B1(_1173_),
    .VDD(VPWR),
    .Y(_0182_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .A2(_1174_));
 sg13g2_nand3b_1 _3113_ (.B(net829),
    .C(net739),
    .Y(_1175_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net830));
 sg13g2_nor3_1 _3114_ (.A(net827),
    .B(net1054),
    .C(_1175_),
    .Y(_1176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3115_ (.A(net397),
    .B(net633),
    .Y(_1177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3116_ (.Y(_1178_),
    .A(net764),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3117_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1178_),
    .Y(_0183_),
    .B1(net398));
 sg13g2_nor2_1 _3118_ (.A(net440),
    .B(net633),
    .Y(_1179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3119_ (.Y(_1180_),
    .A(net762),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3120_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1176_),
    .A2(_1180_),
    .Y(_0184_),
    .B1(net441));
 sg13g2_nor2_1 _3121_ (.A(net325),
    .B(net632),
    .Y(_1181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3122_ (.Y(_1182_),
    .A(net761),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3123_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net632),
    .A2(_1182_),
    .Y(_0185_),
    .B1(_1181_));
 sg13g2_nor2_1 _3124_ (.A(net331),
    .B(net632),
    .Y(_1183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3125_ (.Y(_1184_),
    .A(net760),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3126_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net632),
    .A2(_1184_),
    .Y(_0186_),
    .B1(_1183_));
 sg13g2_nor2_1 _3127_ (.A(net316),
    .B(net632),
    .Y(_1185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3128_ (.Y(_1186_),
    .A(net759),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3129_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net632),
    .A2(_1186_),
    .Y(_0187_),
    .B1(_1185_));
 sg13g2_nor2_1 _3130_ (.A(net358),
    .B(net633),
    .Y(_1187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3131_ (.Y(_1188_),
    .A(\u_usb_cdc.sie_out_data[5] ),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3132_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1188_),
    .Y(_0188_),
    .B1(net359));
 sg13g2_nor2_1 _3133_ (.A(net345),
    .B(net632),
    .Y(_1189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3134_ (.Y(_1190_),
    .A(net758),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3135_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net632),
    .A2(_1190_),
    .Y(_0189_),
    .B1(_1189_));
 sg13g2_nor2_1 _3136_ (.A(net333),
    .B(net633),
    .Y(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3137_ (.Y(_1192_),
    .A(net757),
    .B(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3138_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1192_),
    .Y(_0190_),
    .B1(net334));
 sg13g2_nand2_2 _3139_ (.Y(_1193_),
    .A(net830),
    .B(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3140_ (.A(_1158_),
    .B(_1193_),
    .Y(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3141_ (.Y(_1195_),
    .A(net711),
    .B(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3142_ (.Y(_1196_),
    .A(net172),
    .B(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3143_ (.B1(_1196_),
    .VDD(VPWR),
    .Y(_0191_),
    .VSS(VGND),
    .A1(net723),
    .A2(net605));
 sg13g2_nand2_1 _3144_ (.Y(_1197_),
    .A(net145),
    .B(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3145_ (.B1(_1197_),
    .VDD(VPWR),
    .Y(_0192_),
    .VSS(VGND),
    .A1(net722),
    .A2(net606));
 sg13g2_nor2_1 _3146_ (.A(net761),
    .B(net605),
    .Y(_1198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3147_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1995_),
    .A2(net605),
    .Y(_0193_),
    .B1(_1198_));
 sg13g2_nand2_1 _3148_ (.Y(_1199_),
    .A(net195),
    .B(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3149_ (.B1(_1199_),
    .VDD(VPWR),
    .Y(_0194_),
    .VSS(VGND),
    .A1(net720),
    .A2(net607));
 sg13g2_nor2_1 _3150_ (.A(net759),
    .B(net605),
    .Y(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3151_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1998_),
    .A2(net605),
    .Y(_0195_),
    .B1(_1200_));
 sg13g2_nor2_1 _3152_ (.A(\u_usb_cdc.sie_out_data[5] ),
    .B(net605),
    .Y(_1201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3153_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1999_),
    .A2(net605),
    .Y(_0196_),
    .B1(_1201_));
 sg13g2_nand2_1 _3154_ (.Y(_1202_),
    .A(net160),
    .B(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3155_ (.B1(_1202_),
    .VDD(VPWR),
    .Y(_0197_),
    .VSS(VGND),
    .A1(_1917_),
    .A2(net607));
 sg13g2_nor2_1 _3156_ (.A(net757),
    .B(net606),
    .Y(_1203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3157_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2002_),
    .A2(net605),
    .Y(_0198_),
    .B1(_1203_));
 sg13g2_or3_1 _3158_ (.A(net711),
    .B(_1153_),
    .C(_1158_),
    .X(_1204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3159_ (.Y(_1205_),
    .A(net257),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3160_ (.B1(_1205_),
    .VDD(VPWR),
    .Y(_0199_),
    .VSS(VGND),
    .A1(_1178_),
    .A2(_1204_));
 sg13g2_nand2_1 _3161_ (.Y(_1206_),
    .A(net143),
    .B(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3162_ (.B1(_1206_),
    .VDD(VPWR),
    .Y(_0200_),
    .VSS(VGND),
    .A1(_1180_),
    .A2(net609));
 sg13g2_nand2_1 _3163_ (.Y(_1207_),
    .A(net180),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3164_ (.B1(_1207_),
    .VDD(VPWR),
    .Y(_0201_),
    .VSS(VGND),
    .A1(_1182_),
    .A2(net608));
 sg13g2_nand2_1 _3165_ (.Y(_1208_),
    .A(net125),
    .B(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3166_ (.B1(_1208_),
    .VDD(VPWR),
    .Y(_0202_),
    .VSS(VGND),
    .A1(_1184_),
    .A2(net609));
 sg13g2_nand2_1 _3167_ (.Y(_1209_),
    .A(net185),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3168_ (.B1(_1209_),
    .VDD(VPWR),
    .Y(_0203_),
    .VSS(VGND),
    .A1(_1186_),
    .A2(net608));
 sg13g2_nand2_1 _3169_ (.Y(_1210_),
    .A(net189),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3170_ (.B1(_1210_),
    .VDD(VPWR),
    .Y(_0204_),
    .VSS(VGND),
    .A1(_1188_),
    .A2(net608));
 sg13g2_nand2_1 _3171_ (.Y(_1211_),
    .A(net246),
    .B(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3172_ (.B1(_1211_),
    .VDD(VPWR),
    .Y(_0205_),
    .VSS(VGND),
    .A1(_1190_),
    .A2(net609));
 sg13g2_nand2_1 _3173_ (.Y(_1212_),
    .A(net212),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3174_ (.B1(_1212_),
    .VDD(VPWR),
    .Y(_0206_),
    .VSS(VGND),
    .A1(_1192_),
    .A2(net609));
 sg13g2_nand4_1 _3175_ (.B(net830),
    .C(net827),
    .A(net739),
    .Y(_1213_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1139_));
 sg13g2_nand2_1 _3176_ (.Y(_1214_),
    .A(net214),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3177_ (.B1(_1214_),
    .VDD(VPWR),
    .Y(_0207_),
    .VSS(VGND),
    .A1(net711),
    .A2(_1160_));
 sg13g2_nand2_1 _3178_ (.Y(_1215_),
    .A(net146),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3179_ (.B1(_1215_),
    .VDD(VPWR),
    .Y(_0208_),
    .VSS(VGND),
    .A1(net712),
    .A2(_1162_));
 sg13g2_nand2_1 _3180_ (.Y(_1216_),
    .A(net175),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3181_ (.B1(_1216_),
    .VDD(VPWR),
    .Y(_0209_),
    .VSS(VGND),
    .A1(net712),
    .A2(_1164_));
 sg13g2_nand2_1 _3182_ (.Y(_1217_),
    .A(net127),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3183_ (.B1(_1217_),
    .VDD(VPWR),
    .Y(_0210_),
    .VSS(VGND),
    .A1(net711),
    .A2(_1166_));
 sg13g2_nand2_1 _3184_ (.Y(_1218_),
    .A(net230),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3185_ (.B1(_1218_),
    .VDD(VPWR),
    .Y(_0211_),
    .VSS(VGND),
    .A1(net712),
    .A2(_1168_));
 sg13g2_nand2_1 _3186_ (.Y(_1219_),
    .A(net162),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3187_ (.B1(_1219_),
    .VDD(VPWR),
    .Y(_0212_),
    .VSS(VGND),
    .A1(net712),
    .A2(_1170_));
 sg13g2_nand2_1 _3188_ (.Y(_1220_),
    .A(net234),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3189_ (.B1(_1220_),
    .VDD(VPWR),
    .Y(_0213_),
    .VSS(VGND),
    .A1(net711),
    .A2(_1172_));
 sg13g2_nand2_1 _3190_ (.Y(_1221_),
    .A(net98),
    .B(_1213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3191_ (.B1(_1221_),
    .VDD(VPWR),
    .Y(_0214_),
    .VSS(VGND),
    .A1(net712),
    .A2(_1174_));
 sg13g2_nor3_2 _3192_ (.A(net711),
    .B(net826),
    .C(_1175_),
    .Y(_1222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3193_ (.A(net317),
    .B(net631),
    .Y(_1223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3194_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net723),
    .A2(net631),
    .Y(_0215_),
    .B1(_1223_));
 sg13g2_nor2_1 _3195_ (.A(net342),
    .B(_1222_),
    .Y(_1224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3196_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net722),
    .A2(net631),
    .Y(_0216_),
    .B1(net343));
 sg13g2_nor2_1 _3197_ (.A(net416),
    .B(net630),
    .Y(_1225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3198_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1913_),
    .A2(net630),
    .Y(_0217_),
    .B1(_1225_));
 sg13g2_nor2_1 _3199_ (.A(net347),
    .B(net630),
    .Y(_1226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3200_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net720),
    .A2(net630),
    .Y(_0218_),
    .B1(_1226_));
 sg13g2_nor2_1 _3201_ (.A(net498),
    .B(net630),
    .Y(_1227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3202_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1915_),
    .A2(net630),
    .Y(_0219_),
    .B1(_1227_));
 sg13g2_nor2_1 _3203_ (.A(net402),
    .B(net630),
    .Y(_1228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3204_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1914_),
    .A2(net630),
    .Y(_0220_),
    .B1(_1228_));
 sg13g2_nor2_1 _3205_ (.A(net426),
    .B(net631),
    .Y(_1229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3206_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1917_),
    .A2(net631),
    .Y(_0221_),
    .B1(_1229_));
 sg13g2_nor2_1 _3207_ (.A(net396),
    .B(net631),
    .Y(_1230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3208_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net719),
    .A2(net631),
    .Y(_0222_),
    .B1(_1230_));
 sg13g2_nand3_1 _3209_ (.B(net829),
    .C(net827),
    .A(net831),
    .Y(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3210_ (.Y(_1232_),
    .A(net828),
    .B(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3211_ (.Y(_1233_),
    .A(net224),
    .B(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3212_ (.B1(_1233_),
    .VDD(VPWR),
    .Y(_0223_),
    .VSS(VGND),
    .A1(net723),
    .A2(net604));
 sg13g2_nand2_1 _3213_ (.Y(_1234_),
    .A(net100),
    .B(_1232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3214_ (.B1(net101),
    .VDD(VPWR),
    .Y(_0224_),
    .VSS(VGND),
    .A1(net722),
    .A2(net604));
 sg13g2_nand2_1 _3215_ (.Y(_1235_),
    .A(net276),
    .B(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3216_ (.B1(_1235_),
    .VDD(VPWR),
    .Y(_0225_),
    .VSS(VGND),
    .A1(_1913_),
    .A2(net603));
 sg13g2_nand2_1 _3217_ (.Y(_1236_),
    .A(net211),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3218_ (.B1(_1236_),
    .VDD(VPWR),
    .Y(_0226_),
    .VSS(VGND),
    .A1(net720),
    .A2(net603));
 sg13g2_nand2_1 _3219_ (.Y(_1237_),
    .A(net303),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3220_ (.B1(_1237_),
    .VDD(VPWR),
    .Y(_0227_),
    .VSS(VGND),
    .A1(_1915_),
    .A2(net603));
 sg13g2_nand2_1 _3221_ (.Y(_1238_),
    .A(net323),
    .B(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3222_ (.B1(_1238_),
    .VDD(VPWR),
    .Y(_0228_),
    .VSS(VGND),
    .A1(_1914_),
    .A2(net603));
 sg13g2_nor2_1 _3223_ (.A(net758),
    .B(net603),
    .Y(_1239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3224_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2001_),
    .A2(net603),
    .Y(_0229_),
    .B1(_1239_));
 sg13g2_nand2_1 _3225_ (.Y(_1240_),
    .A(net148),
    .B(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3226_ (.B1(_1240_),
    .VDD(VPWR),
    .Y(_0230_),
    .VSS(VGND),
    .A1(net719),
    .A2(net604));
 sg13g2_nand2_1 _3227_ (.Y(_1241_),
    .A(net152),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3228_ (.B1(_1241_),
    .VDD(VPWR),
    .Y(_0231_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1178_));
 sg13g2_nand2_1 _3229_ (.Y(_1242_),
    .A(net129),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3230_ (.B1(_1242_),
    .VDD(VPWR),
    .Y(_0232_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1180_));
 sg13g2_nand2_1 _3231_ (.Y(_1243_),
    .A(net207),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3232_ (.B1(_1243_),
    .VDD(VPWR),
    .Y(_0233_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1182_));
 sg13g2_nand2_1 _3233_ (.Y(_1244_),
    .A(net191),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3234_ (.B1(_1244_),
    .VDD(VPWR),
    .Y(_0234_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1184_));
 sg13g2_nand2_1 _3235_ (.Y(_1245_),
    .A(net50),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3236_ (.B1(_1245_),
    .VDD(VPWR),
    .Y(_0235_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1186_));
 sg13g2_nand2_1 _3237_ (.Y(_1246_),
    .A(net226),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3238_ (.B1(_1246_),
    .VDD(VPWR),
    .Y(_0236_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1188_));
 sg13g2_nand2_1 _3239_ (.Y(_1247_),
    .A(net166),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3240_ (.B1(_1247_),
    .VDD(VPWR),
    .Y(_0237_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1190_));
 sg13g2_nand2_1 _3241_ (.Y(_1248_),
    .A(net170),
    .B(_1156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3242_ (.B1(_1248_),
    .VDD(VPWR),
    .Y(_0238_),
    .VSS(VGND),
    .A1(_1155_),
    .A2(_1192_));
 sg13g2_nand3_1 _3243_ (.B(net639),
    .C(_0605_),
    .A(net741),
    .Y(_1249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3244_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1250_),
    .B(_1231_),
    .A(_1981_));
 sg13g2_nand2b_1 _3245_ (.Y(_1251_),
    .B(_1250_),
    .A_N(_1154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3246_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1981_),
    .A2(_1231_),
    .Y(_1252_),
    .B1(_1251_));
 sg13g2_xnor2_1 _3247_ (.Y(_1253_),
    .A(_1983_),
    .B(_1252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3248_ (.Y(_1254_),
    .A(_1153_),
    .B(_1193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3249_ (.B(_1254_),
    .A(net814),
    .X(_1255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3250_ (.Y(_1256_),
    .A(net827),
    .B(_1193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3251_ (.Y(_1257_),
    .A(net813),
    .B(_1256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3252_ (.B(_1255_),
    .C(_1257_),
    .A(_1250_),
    .Y(_1258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3253_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net826),
    .A2(_1154_),
    .Y(_1259_),
    .B1(net831));
 sg13g2_inv_1 _3254_ (.VDD(VPWR),
    .Y(_1260_),
    .A(_1259_),
    .VSS(VGND));
 sg13g2_xor2_1 _3255_ (.B(_1259_),
    .A(net820),
    .X(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3256_ (.A(_1253_),
    .B(_1258_),
    .C(_1261_),
    .Y(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3257_ (.B1(_0714_),
    .VDD(VPWR),
    .Y(_1263_),
    .VSS(VGND),
    .A1(net770),
    .A2(_1262_));
 sg13g2_nand2b_2 _3258_ (.Y(_1264_),
    .B(_1263_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1249_));
 sg13g2_nor2_1 _3259_ (.A(net770),
    .B(net830),
    .Y(_1265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3260_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net771),
    .A2(_1984_),
    .Y(_1266_),
    .B1(_1265_));
 sg13g2_nor3_1 _3261_ (.A(net755),
    .B(_0601_),
    .C(_1266_),
    .Y(_1267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3262_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1260_),
    .C1(_1267_),
    .B1(_0714_),
    .A1(net755),
    .Y(_1268_),
    .A2(_1984_));
 sg13g2_mux2_1 _3263_ (.A0(_1268_),
    .A1(net830),
    .S(_1264_),
    .X(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3264_ (.A0(net829),
    .A1(net935),
    .S(net770),
    .X(_1269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3265_ (.B(_1153_),
    .C(_1193_),
    .A(_0714_),
    .Y(_1270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3266_ (.Y(_1271_),
    .B1(_0604_),
    .B2(_1269_),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .A1(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3267_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1270_),
    .A2(_1271_),
    .Y(_1272_),
    .B1(_1264_));
 sg13g2_a21o_1 _3268_ (.A2(_1264_),
    .A1(net892),
    .B1(_1272_),
    .X(_0240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3269_ (.Y(_1273_),
    .A(net770),
    .B(net940),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3270_ (.B1(_1273_),
    .VDD(VPWR),
    .Y(_1274_),
    .VSS(VGND),
    .A1(net770),
    .A2(net711));
 sg13g2_nand2_1 _3271_ (.Y(_1275_),
    .A(_0714_),
    .B(_1256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3272_ (.Y(_1276_),
    .B1(_0604_),
    .B2(_1274_),
    .A2(net940),
    .A1(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1275_),
    .A2(_1276_),
    .Y(_1277_),
    .B1(_1264_));
 sg13g2_a21o_1 _3274_ (.A2(_1264_),
    .A1(net828),
    .B1(_1277_),
    .X(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3275_ (.Y(_1278_),
    .A(_0714_),
    .B(_1252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3276_ (.Y(_1279_),
    .A(net770),
    .B(net951),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3277_ (.B1(_1279_),
    .VDD(VPWR),
    .Y(_1280_),
    .VSS(VGND),
    .A1(net770),
    .A2(_1981_));
 sg13g2_a22oi_1 _3278_ (.Y(_1281_),
    .B1(_0604_),
    .B2(_1280_),
    .A2(net951),
    .A1(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3279_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1278_),
    .A2(_1281_),
    .Y(_1282_),
    .B1(_1264_));
 sg13g2_a21o_1 _3280_ (.A2(_1264_),
    .A1(net826),
    .B1(_1282_),
    .X(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3281_ (.A(_0936_),
    .B_N(_0937_),
    .Y(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3282_ (.Y(_1284_),
    .B(_0937_),
    .A_N(_0936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3283_ (.S0(net824),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .S1(net816),
    .X(_1285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3284_ (.Y(_1286_),
    .A(net816),
    .B(_1982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3285_ (.A(net816),
    .B(net812),
    .Y(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3286_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1288_),
    .B(net813),
    .A(net814));
 sg13g2_mux2_1 _3287_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .S(net824),
    .X(_1289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3288_ (.A(net823),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .Y(_1290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3289_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .B_N(net821),
    .Y(_1291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3290_ (.A(_1286_),
    .B(_1290_),
    .C(_1291_),
    .Y(_1292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3291_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1289_),
    .C1(_1292_),
    .B1(_1287_),
    .A1(net812),
    .Y(_1293_),
    .A2(_1285_));
 sg13g2_nor3_2 _3292_ (.A(net819),
    .B(_1983_),
    .C(_1288_),
    .Y(_1294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3293_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net152),
    .A2(net629),
    .Y(_1295_),
    .B1(net617));
 sg13g2_o21ai_1 _3294_ (.B1(_1295_),
    .VDD(VPWR),
    .Y(_1296_),
    .VSS(VGND),
    .A1(net965),
    .A2(_1293_));
 sg13g2_o21ai_1 _3295_ (.B1(_1296_),
    .VDD(VPWR),
    .Y(_1297_),
    .VSS(VGND),
    .A1(net985),
    .A2(_1283_));
 sg13g2_inv_1 _3296_ (.VDD(VPWR),
    .Y(_0243_),
    .A(_1297_),
    .VSS(VGND));
 sg13g2_mux4_1 _3297_ (.S0(net825),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .S1(net817),
    .X(_1298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3298_ (.Y(_1299_),
    .B(net822),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3299_ (.B1(_1299_),
    .VDD(VPWR),
    .Y(_1300_),
    .VSS(VGND),
    .A1(net822),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ));
 sg13g2_mux2_1 _3300_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .S(net824),
    .X(_1301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3301_ (.Y(_1302_),
    .B1(_1301_),
    .B2(_1287_),
    .A2(_1298_),
    .A1(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3302_ (.B1(_1302_),
    .VDD(VPWR),
    .Y(_1303_),
    .VSS(VGND),
    .A1(_1286_),
    .A2(_1300_));
 sg13g2_a221oi_1 _3303_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1983_),
    .C1(net616),
    .B1(_1303_),
    .A1(net129),
    .Y(_1304_),
    .A2(net629));
 sg13g2_a21oi_1 _3304_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2008_),
    .A2(net616),
    .Y(_0244_),
    .B1(_1304_));
 sg13g2_mux4_1 _3305_ (.S0(net821),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .S1(net816),
    .X(_1305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3306_ (.Y(_1306_),
    .B(net822),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3307_ (.B1(_1306_),
    .VDD(VPWR),
    .Y(_1307_),
    .VSS(VGND),
    .A1(net822),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ));
 sg13g2_or2_1 _3308_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1308_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[18] ),
    .A(net823));
 sg13g2_a21oi_1 _3309_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net821),
    .A2(_1995_),
    .Y(_1309_),
    .B1(_1286_));
 sg13g2_a22oi_1 _3310_ (.Y(_1310_),
    .B1(_1308_),
    .B2(_1309_),
    .A2(_1305_),
    .A1(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3311_ (.B1(_1310_),
    .VDD(VPWR),
    .Y(_1311_),
    .VSS(VGND),
    .A1(_1288_),
    .A2(_1307_));
 sg13g2_a221oi_1 _3312_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1983_),
    .C1(net616),
    .B1(_1311_),
    .A1(net207),
    .Y(_1312_),
    .A2(net629));
 sg13g2_a21oi_1 _3313_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2009_),
    .A2(net616),
    .Y(_0245_),
    .B1(_1312_));
 sg13g2_nor2_1 _3314_ (.A(net445),
    .B(_1283_),
    .Y(_1313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3315_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net818),
    .A2(_1996_),
    .Y(_1314_),
    .B1(net814));
 sg13g2_o21ai_1 _3316_ (.B1(_1314_),
    .VDD(VPWR),
    .Y(_1315_),
    .VSS(VGND),
    .A1(net818),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[3] ));
 sg13g2_mux2_1 _3317_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .S(net818),
    .X(_1316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3318_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net815),
    .A2(_1316_),
    .Y(_1317_),
    .B1(net812));
 sg13g2_a21oi_1 _3319_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net818),
    .A2(_1997_),
    .Y(_1318_),
    .B1(net815));
 sg13g2_o21ai_1 _3320_ (.B1(_1318_),
    .VDD(VPWR),
    .Y(_1319_),
    .VSS(VGND),
    .A1(net818),
    .A2(net125));
 sg13g2_mux2_1 _3321_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[51] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[59] ),
    .S(net821),
    .X(_1320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3322_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net816),
    .A2(_1320_),
    .Y(_1321_),
    .B1(_1982_));
 sg13g2_a22oi_1 _3323_ (.Y(_1322_),
    .B1(_1319_),
    .B2(_1321_),
    .A2(_1317_),
    .A1(_1315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3324_ (.Y(_1323_),
    .B1(_1322_),
    .B2(_1983_),
    .A2(net629),
    .A1(net191),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3325_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1283_),
    .A2(_1323_),
    .Y(_0246_),
    .B1(net446));
 sg13g2_mux4_1 _3326_ (.S0(net823),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .S1(net816),
    .X(_1324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3327_ (.Y(_1325_),
    .B(net823),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3328_ (.B1(_1325_),
    .VDD(VPWR),
    .Y(_1326_),
    .VSS(VGND),
    .A1(net823),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ));
 sg13g2_or2_1 _3329_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1327_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .A(net823));
 sg13g2_a21oi_1 _3330_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net821),
    .A2(_1998_),
    .Y(_1328_),
    .B1(_1286_));
 sg13g2_a22oi_1 _3331_ (.Y(_1329_),
    .B1(_1327_),
    .B2(_1328_),
    .A2(_1324_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3332_ (.B1(_1329_),
    .VDD(VPWR),
    .Y(_1330_),
    .VSS(VGND),
    .A1(_1288_),
    .A2(_1326_));
 sg13g2_a221oi_1 _3333_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1983_),
    .C1(net616),
    .B1(_1330_),
    .A1(net50),
    .Y(_1331_),
    .A2(net629));
 sg13g2_a21oi_1 _3334_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2010_),
    .A2(net616),
    .Y(_0247_),
    .B1(net51));
 sg13g2_mux4_1 _3335_ (.S0(net821),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .S1(net816),
    .X(_1332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3336_ (.Y(_1333_),
    .B(net825),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3337_ (.B1(_1333_),
    .VDD(VPWR),
    .Y(_1334_),
    .VSS(VGND),
    .A1(net822),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ));
 sg13g2_or2_1 _3338_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1335_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .A(net823));
 sg13g2_a21oi_1 _3339_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net822),
    .A2(_1999_),
    .Y(_1336_),
    .B1(_1286_));
 sg13g2_a22oi_1 _3340_ (.Y(_1337_),
    .B1(_1335_),
    .B2(_1336_),
    .A2(_1332_),
    .A1(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3341_ (.B1(_1337_),
    .VDD(VPWR),
    .Y(_1338_),
    .VSS(VGND),
    .A1(_1288_),
    .A2(_1334_));
 sg13g2_a221oi_1 _3342_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1983_),
    .C1(net617),
    .B1(_1338_),
    .A1(net226),
    .Y(_1339_),
    .A2(_1294_));
 sg13g2_a21oi_1 _3343_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2011_),
    .A2(net616),
    .Y(_0248_),
    .B1(_1339_));
 sg13g2_a21oi_1 _3344_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net819),
    .A2(_2000_),
    .Y(_1340_),
    .B1(net815));
 sg13g2_o21ai_1 _3345_ (.B1(_1340_),
    .VDD(VPWR),
    .Y(_1341_),
    .VSS(VGND),
    .A1(net819),
    .A2(net255));
 sg13g2_mux2_1 _3346_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .S(net818),
    .X(_1342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3347_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net815),
    .A2(_1342_),
    .Y(_1343_),
    .B1(net813));
 sg13g2_nand2b_1 _3348_ (.Y(_1344_),
    .B(net818),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3349_ (.B1(_1344_),
    .VDD(VPWR),
    .Y(_1345_),
    .VSS(VGND),
    .A1(net818),
    .A2(net246));
 sg13g2_o21ai_1 _3350_ (.B1(net816),
    .VDD(VPWR),
    .Y(_1346_),
    .VSS(VGND),
    .A1(net821),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[54] ));
 sg13g2_a21oi_1 _3351_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net821),
    .A2(_2001_),
    .Y(_1347_),
    .B1(_1346_));
 sg13g2_o21ai_1 _3352_ (.B1(net813),
    .VDD(VPWR),
    .Y(_1348_),
    .VSS(VGND),
    .A1(net814),
    .A2(_1345_));
 sg13g2_a21oi_1 _3353_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1341_),
    .A2(_1343_),
    .Y(_1349_),
    .B1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ));
 sg13g2_o21ai_1 _3354_ (.B1(_1349_),
    .VDD(VPWR),
    .Y(_1350_),
    .VSS(VGND),
    .A1(_1347_),
    .A2(_1348_));
 sg13g2_a21oi_1 _3355_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net166),
    .A2(net629),
    .Y(_1351_),
    .B1(net617));
 sg13g2_a22oi_1 _3356_ (.Y(_0249_),
    .B1(_1350_),
    .B2(_1351_),
    .A2(net616),
    .A1(_2012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3357_ (.S0(net824),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .S1(net817),
    .X(_1352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3358_ (.Y(_1353_),
    .B(net824),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3359_ (.B1(_1353_),
    .VDD(VPWR),
    .Y(_1354_),
    .VSS(VGND),
    .A1(net824),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ));
 sg13g2_or2_1 _3360_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1355_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[23] ),
    .A(net824));
 sg13g2_a21oi_1 _3361_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net824),
    .A2(_2002_),
    .Y(_1356_),
    .B1(_1286_));
 sg13g2_a22oi_1 _3362_ (.Y(_1357_),
    .B1(_1355_),
    .B2(_1356_),
    .A2(_1352_),
    .A1(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3363_ (.B1(_1357_),
    .VDD(VPWR),
    .Y(_1358_),
    .VSS(VGND),
    .A1(_1288_),
    .A2(_1354_));
 sg13g2_a221oi_1 _3364_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1983_),
    .C1(net617),
    .B1(_1358_),
    .A1(net170),
    .Y(_1359_),
    .A2(_1294_));
 sg13g2_a21oi_1 _3365_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2013_),
    .A2(net617),
    .Y(_0250_),
    .B1(_1359_));
 sg13g2_nor3_2 _3366_ (.A(net755),
    .B(_0601_),
    .C(_1249_),
    .Y(_1360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3367_ (.Y(_1361_),
    .A(_1266_),
    .B(_1360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3368_ (.B1(_1361_),
    .VDD(VPWR),
    .Y(_0251_),
    .VSS(VGND),
    .A1(_1984_),
    .A2(_1360_));
 sg13g2_mux2_1 _3369_ (.A0(net935),
    .A1(_1269_),
    .S(_1360_),
    .X(_0252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3370_ (.A0(net940),
    .A1(_1274_),
    .S(_1360_),
    .X(_0253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3371_ (.A0(net951),
    .A1(_1280_),
    .S(_1360_),
    .X(_0254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3372_ (.Y(_1362_),
    .A(net820),
    .B(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3373_ (.A(net629),
    .B(_1362_),
    .Y(_0255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3374_ (.B(net814),
    .C(_1283_),
    .A(net820),
    .Y(_1363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3375_ (.A2(_1283_),
    .A1(net820),
    .B1(net814),
    .X(_1364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3376_ (.A(_1363_),
    .B(_1364_),
    .X(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3377_ (.Y(_0257_),
    .A(net813),
    .B(_1363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3378_ (.B(net814),
    .C(net813),
    .A(net820),
    .Y(_1365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3379_ (.A(net629),
    .B_N(_1365_),
    .Y(_1366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3380_ (.B1(net965),
    .VDD(VPWR),
    .Y(_1367_),
    .VSS(VGND),
    .A1(net617),
    .A2(_1366_));
 sg13g2_or2_1 _3381_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1368_),
    .B(_1365_),
    .A(net617));
 sg13g2_o21ai_1 _3382_ (.B1(_1367_),
    .VDD(VPWR),
    .Y(_0258_),
    .VSS(VGND),
    .A1(net965),
    .A2(_1368_));
 sg13g2_nand2_2 _3383_ (.Y(_1369_),
    .A(_1128_),
    .B(_1134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3384_ (.B(net931),
    .C(net639),
    .A(net1034),
    .Y(_1370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3385_ (.A(net809),
    .B(net801),
    .C(net797),
    .Y(_1371_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1924_));
 sg13g2_a21o_1 _3386_ (.A2(net639),
    .A1(\u_usb_cdc.sie_in_req ),
    .B1(_1371_),
    .X(_1372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3387_ (.B1(_1370_),
    .VDD(VPWR),
    .Y(_1373_),
    .VSS(VGND),
    .A1(net809),
    .A2(_1372_));
 sg13g2_mux2_1 _3388_ (.A0(_1373_),
    .A1(net811),
    .S(_1369_),
    .X(_0259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3389_ (.Y(_1374_),
    .A(net809),
    .B(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3390_ (.Y(_1375_),
    .A(_1133_),
    .B(_1374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3391_ (.B1(_1375_),
    .VDD(VPWR),
    .Y(_1376_),
    .VSS(VGND),
    .A1(net575),
    .A2(_1133_));
 sg13g2_nand2_1 _3392_ (.Y(_1377_),
    .A(net802),
    .B(_1369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3393_ (.B1(net1015),
    .VDD(VPWR),
    .Y(_0260_),
    .VSS(VGND),
    .A1(_1369_),
    .A2(_1376_));
 sg13g2_nor2_1 _3394_ (.A(net419),
    .B(_1133_),
    .Y(_1378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3395_ (.B(net802),
    .C(net797),
    .A(net809),
    .Y(_1379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3396_ (.A2(net802),
    .A1(net809),
    .B1(net797),
    .X(_1380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3397_ (.Y(_1381_),
    .A(_1379_),
    .B(_1380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3398_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1133_),
    .A2(_1381_),
    .Y(_1382_),
    .B1(_1378_));
 sg13g2_nor2_1 _3399_ (.A(_1369_),
    .B(_1382_),
    .Y(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3400_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1923_),
    .A2(_1369_),
    .Y(_0261_),
    .B1(_1383_));
 sg13g2_nand3_1 _3401_ (.B(net363),
    .C(net639),
    .A(\u_usb_cdc.sie_in_req ),
    .Y(_1384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3402_ (.Y(_1385_),
    .A(_1924_),
    .B(_1379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3403_ (.B1(_1384_),
    .VDD(VPWR),
    .Y(_1386_),
    .VSS(VGND),
    .A1(_1372_),
    .A2(_1385_));
 sg13g2_mux2_1 _3404_ (.A0(_1386_),
    .A1(net980),
    .S(_1369_),
    .X(_0262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3405_ (.A(net624),
    .B(_0671_),
    .Y(_1387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3406_ (.A(_0611_),
    .B(_0616_),
    .C(_0644_),
    .Y(_1388_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0665_));
 sg13g2_nand2_2 _3407_ (.Y(_1389_),
    .A(net743),
    .B(_1388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3408_ (.A(_1387_),
    .B(_1389_),
    .Y(_1390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3409_ (.A(net418),
    .B(net578),
    .Y(_1391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3410_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net724),
    .A2(net578),
    .Y(_0263_),
    .B1(_1391_));
 sg13g2_nor2_1 _3411_ (.A(net871),
    .B(net578),
    .Y(_1392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3412_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net721),
    .A2(_1390_),
    .Y(_0264_),
    .B1(_1392_));
 sg13g2_nor2_1 _3413_ (.A(net545),
    .B(net578),
    .Y(_1393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3414_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1913_),
    .A2(net578),
    .Y(_0265_),
    .B1(_1393_));
 sg13g2_nor2_1 _3415_ (.A(net500),
    .B(net578),
    .Y(_1394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3416_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net720),
    .A2(net578),
    .Y(_0266_),
    .B1(_1394_));
 sg13g2_nor2_1 _3417_ (.A(net901),
    .B(net578),
    .Y(_1395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3418_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net719),
    .A2(_1390_),
    .Y(_0267_),
    .B1(_1395_));
 sg13g2_nor2b_1 _3419_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .B_N(net849),
    .Y(_1396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3420_ (.A(_0588_),
    .B(_0623_),
    .C(_1396_),
    .Y(_1397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3421_ (.A0(net868),
    .A1(net499),
    .S(_1397_),
    .X(_0268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3422_ (.A0(net905),
    .A1(net485),
    .S(_1397_),
    .X(_0269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3423_ (.A0(net861),
    .A1(net428),
    .S(_1397_),
    .X(_0270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3424_ (.A0(net923),
    .A1(net559),
    .S(_1397_),
    .X(_0271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3425_ (.A0(net897),
    .A1(net566),
    .S(_1397_),
    .X(_0272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3426_ (.A0(net878),
    .A1(net473),
    .S(_1397_),
    .X(_0273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3427_ (.A0(net900),
    .A1(net435),
    .S(_1397_),
    .X(_0274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3428_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net850),
    .A2(_0601_),
    .Y(_1398_),
    .B1(net715));
 sg13g2_nor3_1 _3429_ (.A(\u_usb_cdc.sie_out_data[7] ),
    .B(_1941_),
    .C(_0640_),
    .Y(_1399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3430_ (.A(_1398_),
    .B(_1399_),
    .Y(_1400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3431_ (.A(_1400_),
    .B_N(_1388_),
    .Y(_1401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3432_ (.A(net499),
    .B(net582),
    .Y(_1402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3433_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net724),
    .A2(net582),
    .Y(_0275_),
    .B1(_1402_));
 sg13g2_nor2_1 _3434_ (.A(net485),
    .B(net582),
    .Y(_1403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3435_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net721),
    .A2(net582),
    .Y(_0276_),
    .B1(_1403_));
 sg13g2_nor2_1 _3436_ (.A(net428),
    .B(net581),
    .Y(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3437_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1913_),
    .A2(net581),
    .Y(_0277_),
    .B1(_1404_));
 sg13g2_nor2_1 _3438_ (.A(net559),
    .B(net582),
    .Y(_1405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net720),
    .A2(net582),
    .Y(_0278_),
    .B1(_1405_));
 sg13g2_nor2_1 _3440_ (.A(net566),
    .B(net581),
    .Y(_1406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3441_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1915_),
    .A2(net581),
    .Y(_0279_),
    .B1(_1406_));
 sg13g2_nor2_1 _3442_ (.A(net473),
    .B(net581),
    .Y(_1407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3443_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1914_),
    .A2(net581),
    .Y(_0280_),
    .B1(_1407_));
 sg13g2_nor2_1 _3444_ (.A(net435),
    .B(net581),
    .Y(_1408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3445_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1917_),
    .A2(net581),
    .Y(_0281_),
    .B1(_1408_));
 sg13g2_nor3_1 _3446_ (.A(_1940_),
    .B(_0640_),
    .C(_0693_),
    .Y(_1409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3447_ (.B1(_1388_),
    .VDD(VPWR),
    .Y(_1410_),
    .VSS(VGND),
    .A1(_1398_),
    .A2(_1409_));
 sg13g2_mux2_1 _3448_ (.A0(net623),
    .A1(net489),
    .S(_1410_),
    .X(_0282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3449_ (.Y(_0283_),
    .B(_1410_),
    .A_N(net179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3450_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0634_),
    .A2(_0685_),
    .Y(_1411_),
    .B1(net624));
 sg13g2_nor2_2 _3451_ (.A(_1389_),
    .B(_1411_),
    .Y(_1412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3452_ (.A(net880),
    .B(_1412_),
    .Y(_1413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3453_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net724),
    .A2(_1412_),
    .Y(_0284_),
    .B1(_1413_));
 sg13g2_nor2_1 _3454_ (.A(net953),
    .B(_1412_),
    .Y(_1414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3455_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net722),
    .A2(_1412_),
    .Y(_0285_),
    .B1(_1414_));
 sg13g2_nor2_1 _3456_ (.A(net492),
    .B(_1412_),
    .Y(_1415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3457_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1914_),
    .A2(_1412_),
    .Y(_0286_),
    .B1(_1415_));
 sg13g2_nor2_1 _3458_ (.A(net794),
    .B(_1412_),
    .Y(_1416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3459_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net719),
    .A2(_1412_),
    .Y(_0287_),
    .B1(_1416_));
 sg13g2_nor3_1 _3460_ (.A(_0661_),
    .B(net622),
    .C(_0751_),
    .Y(_1417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3461_ (.A(net624),
    .B(_0648_),
    .C(_1417_),
    .Y(_1418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3462_ (.A(_1389_),
    .B(_1418_),
    .Y(_1419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3463_ (.A(net881),
    .B(net576),
    .Y(_1420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3464_ (.B1(_0661_),
    .VDD(VPWR),
    .Y(_1421_),
    .VSS(VGND),
    .A1(net719),
    .A2(_0751_));
 sg13g2_nor2_1 _3465_ (.A(net763),
    .B(_1421_),
    .Y(_1422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3466_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net576),
    .A2(_1422_),
    .Y(_0288_),
    .B1(_1420_));
 sg13g2_nor2_1 _3467_ (.A(net926),
    .B(net576),
    .Y(_1423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3468_ (.A(\u_usb_cdc.sie_out_data[1] ),
    .B(_1421_),
    .Y(_1424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3469_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net576),
    .A2(_1424_),
    .Y(_0289_),
    .B1(_1423_));
 sg13g2_nor2_1 _3470_ (.A(net864),
    .B(net576),
    .Y(_1425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3471_ (.A(\u_usb_cdc.sie_out_data[2] ),
    .B(_1421_),
    .Y(_1426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3472_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net576),
    .A2(_1426_),
    .Y(_0290_),
    .B1(_1425_));
 sg13g2_nor2_1 _3473_ (.A(net898),
    .B(net576),
    .Y(_1427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3474_ (.A(net760),
    .B(_1421_),
    .Y(_1428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3475_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net576),
    .A2(_1428_),
    .Y(_0291_),
    .B1(_1427_));
 sg13g2_nor2_1 _3476_ (.A(net922),
    .B(net577),
    .Y(_1429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3477_ (.A(net298),
    .B(_1421_),
    .Y(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3478_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_1430_),
    .Y(_0292_),
    .B1(_1429_));
 sg13g2_nor2_1 _3479_ (.A(net908),
    .B(net577),
    .Y(_1431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3480_ (.A(\u_usb_cdc.sie_out_data[5] ),
    .B(_1421_),
    .Y(_1432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3481_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_1432_),
    .Y(_0293_),
    .B1(_1431_));
 sg13g2_nor2_1 _3482_ (.A(net564),
    .B(net577),
    .Y(_1433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3483_ (.A(\u_usb_cdc.sie_out_data[6] ),
    .B(_1421_),
    .Y(_1434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3484_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_1434_),
    .Y(_0294_),
    .B1(_1433_));
 sg13g2_a21oi_1 _3485_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0549_),
    .A2(_0624_),
    .Y(_1435_),
    .B1(_1929_));
 sg13g2_nor2_1 _3486_ (.A(net849),
    .B(_1435_),
    .Y(_1436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3487_ (.B1(_0619_),
    .VDD(VPWR),
    .Y(_1437_),
    .VSS(VGND),
    .A1(_0621_),
    .A2(_1436_));
 sg13g2_o21ai_1 _3488_ (.B1(_1929_),
    .VDD(VPWR),
    .Y(_1438_),
    .VSS(VGND),
    .A1(_0551_),
    .A2(_0602_));
 sg13g2_nand3_1 _3489_ (.B(_1436_),
    .C(_1438_),
    .A(net588),
    .Y(_1439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3490_ (.Y(_1440_),
    .A(net793),
    .B(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3491_ (.B1(_1440_),
    .VDD(VPWR),
    .Y(_0295_),
    .VSS(VGND),
    .A1(net793),
    .A2(_1439_));
 sg13g2_nor2_2 _3492_ (.A(_0540_),
    .B(_0668_),
    .Y(_1441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3493_ (.A(_1439_),
    .B_N(_1441_),
    .Y(_1442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3494_ (.A2(_1437_),
    .A1(net789),
    .B1(_1442_),
    .X(_0296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3495_ (.Y(_1443_),
    .A(net786),
    .B(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3496_ (.Y(_1444_),
    .A(net786),
    .B(_0540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3497_ (.B1(_1443_),
    .VDD(VPWR),
    .Y(_0297_),
    .VSS(VGND),
    .A1(_1439_),
    .A2(_1444_));
 sg13g2_nand2_1 _3498_ (.Y(_1445_),
    .A(net781),
    .B(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3499_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1446_),
    .B(_0655_),
    .A(_0541_));
 sg13g2_nand2_1 _3500_ (.Y(_1447_),
    .A(_0653_),
    .B(_1446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3501_ (.B1(_1445_),
    .VDD(VPWR),
    .Y(_0298_),
    .VSS(VGND),
    .A1(_1439_),
    .A2(_1447_));
 sg13g2_nand2_1 _3502_ (.Y(_1448_),
    .A(net778),
    .B(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3503_ (.B(net781),
    .C(net776),
    .A(net785),
    .Y(_1449_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0540_));
 sg13g2_xor2_1 _3504_ (.B(_1446_),
    .A(net778),
    .X(_1450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3505_ (.B1(_1448_),
    .VDD(VPWR),
    .Y(_0299_),
    .VSS(VGND),
    .A1(_1439_),
    .A2(_1450_));
 sg13g2_nand2_1 _3506_ (.Y(_1451_),
    .A(net774),
    .B(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3507_ (.Y(_1452_),
    .A(net778),
    .B(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3508_ (.A(_1446_),
    .B(_1452_),
    .Y(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3509_ (.B(_1449_),
    .A(net774),
    .X(_1454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3510_ (.B1(_1451_),
    .VDD(VPWR),
    .Y(_0300_),
    .VSS(VGND),
    .A1(_1439_),
    .A2(_1454_));
 sg13g2_nand2_1 _3511_ (.Y(_1455_),
    .A(net562),
    .B(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3512_ (.Y(_1456_),
    .A(net562),
    .B(_1453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3513_ (.B1(_1455_),
    .VDD(VPWR),
    .Y(_0301_),
    .VSS(VGND),
    .A1(_1439_),
    .A2(_1456_));
 sg13g2_nand2b_1 _3514_ (.Y(_1457_),
    .B(_1249_),
    .A_N(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3515_ (.A(_1264_),
    .B(_1457_),
    .X(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3516_ (.A(net993),
    .B(net586),
    .Y(_1458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3517_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net719),
    .A2(net586),
    .Y(_0303_),
    .B1(_1458_));
 sg13g2_mux2_1 _3518_ (.A0(net995),
    .A1(net767),
    .S(net587),
    .X(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3519_ (.A0(net972),
    .A1(net766),
    .S(net587),
    .X(_0305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3520_ (.A0(net971),
    .A1(net765),
    .S(net587),
    .X(_0306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3521_ (.A(net449),
    .B(net586),
    .Y(_1459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3522_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net721),
    .A2(net586),
    .Y(_0307_),
    .B1(_1459_));
 sg13g2_nor2_1 _3523_ (.A(net385),
    .B(net585),
    .Y(_1460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3524_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1913_),
    .A2(net585),
    .Y(_0308_),
    .B1(_1460_));
 sg13g2_nor2_1 _3525_ (.A(net448),
    .B(net585),
    .Y(_1461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3526_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net720),
    .A2(net585),
    .Y(_0309_),
    .B1(_1461_));
 sg13g2_nor2_1 _3527_ (.A(net408),
    .B(net585),
    .Y(_1462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3528_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1915_),
    .A2(net585),
    .Y(_0310_),
    .B1(_1462_));
 sg13g2_nor2_1 _3529_ (.A(net381),
    .B(net586),
    .Y(_1463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3530_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1914_),
    .A2(net586),
    .Y(_0311_),
    .B1(_1463_));
 sg13g2_nor2_1 _3531_ (.A(net409),
    .B(net585),
    .Y(_1464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3532_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1917_),
    .A2(net585),
    .Y(_0312_),
    .B1(_1464_));
 sg13g2_a21oi_1 _3533_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1940_),
    .A2(_1396_),
    .Y(_1465_),
    .B1(_0588_));
 sg13g2_a22oi_1 _3534_ (.Y(_1466_),
    .B1(_0619_),
    .B2(_1465_),
    .A2(\u_usb_cdc.bus_reset ),
    .A1(net742),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3535_ (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[2] ),
    .B(\u_usb_cdc.u_ctrl_endp.addr_dd[5] ),
    .C(\u_usb_cdc.u_ctrl_endp.addr_dd[4] ),
    .D(\u_usb_cdc.u_ctrl_endp.addr_dd[6] ),
    .Y(_1467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3536_ (.A(net851),
    .B(\u_usb_cdc.u_ctrl_endp.addr_dd[1] ),
    .C(\u_usb_cdc.u_ctrl_endp.addr_dd[0] ),
    .D(\u_usb_cdc.u_ctrl_endp.addr_dd[3] ),
    .Y(_1468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3537_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net917),
    .Y(_1469_),
    .A2(_1468_),
    .A1(_1467_));
 sg13g2_o21ai_1 _3538_ (.B1(_1469_),
    .VDD(VPWR),
    .Y(_1470_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1940_));
 sg13g2_mux2_1 _3539_ (.A0(_1470_),
    .A1(net955),
    .S(_1466_),
    .X(_0313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3540_ (.Y(_1471_),
    .A(net413),
    .B(_1466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3541_ (.B1(_1469_),
    .VDD(VPWR),
    .Y(_1472_),
    .VSS(VGND),
    .A1(_1940_),
    .A2(net179));
 sg13g2_o21ai_1 _3542_ (.B1(net414),
    .VDD(VPWR),
    .Y(_0314_),
    .VSS(VGND),
    .A1(_1466_),
    .A2(_1472_));
 sg13g2_nor4_1 _3543_ (.A(net753),
    .B(net717),
    .C(_0436_),
    .D(_0841_),
    .Y(_1473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3544_ (.A2(net717),
    .A1(net1034),
    .B1(_1473_),
    .X(_0315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3545_ (.A(net844),
    .B(_0951_),
    .Y(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3546_ (.Y(_1475_),
    .A(_1972_),
    .B(_0950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3547_ (.B1(net745),
    .VDD(VPWR),
    .Y(_1476_),
    .VSS(VGND),
    .A1(_0603_),
    .A2(_1475_));
 sg13g2_nand3_1 _3548_ (.B(_0603_),
    .C(_1474_),
    .A(net745),
    .Y(_1477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3549_ (.Y(_1478_),
    .A(net354),
    .B(_1476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3550_ (.B1(_1478_),
    .VDD(VPWR),
    .Y(_0316_),
    .VSS(VGND),
    .A1(net354),
    .A2(_1477_));
 sg13g2_nand2_1 _3551_ (.Y(_1479_),
    .A(net430),
    .B(_1476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3552_ (.Y(_1480_),
    .A(net430),
    .B(net354),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3553_ (.B1(net431),
    .VDD(VPWR),
    .Y(_0317_),
    .VSS(VGND),
    .A1(_1477_),
    .A2(_1480_));
 sg13g2_nand3_1 _3554_ (.B(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .C(net745),
    .A(\u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .Y(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3555_ (.Y(_0318_),
    .B1(_1481_),
    .B2(_1930_),
    .A2(_1475_),
    .A1(net746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3556_ (.Y(_1482_),
    .A(net327),
    .B(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3557_ (.B1(_1482_),
    .VDD(VPWR),
    .Y(_0319_),
    .VSS(VGND),
    .A1(net327),
    .A2(_0867_));
 sg13g2_nand2_1 _3558_ (.Y(_1483_),
    .A(net376),
    .B(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3559_ (.Y(_1484_),
    .A(net376),
    .B(net327),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3560_ (.B1(_1483_),
    .VDD(VPWR),
    .Y(_0320_),
    .VSS(VGND),
    .A1(_0867_),
    .A2(_1484_));
 sg13g2_nand2_1 _3561_ (.Y(_1485_),
    .A(net321),
    .B(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3562_ (.A2(\u_usb_cdc.u_sie.in_byte_q[0] ),
    .A1(\u_usb_cdc.u_sie.in_byte_q[1] ),
    .B1(net321),
    .X(_1486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3563_ (.Y(_1487_),
    .A(_0584_),
    .B(_1486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3564_ (.B1(_1485_),
    .VDD(VPWR),
    .Y(_0321_),
    .VSS(VGND),
    .A1(_0867_),
    .A2(_1487_));
 sg13g2_nand2_1 _3565_ (.Y(_1488_),
    .A(net400),
    .B(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3566_ (.B(_0584_),
    .A(net400),
    .X(_1489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3567_ (.B1(_1488_),
    .VDD(VPWR),
    .Y(_0322_),
    .VSS(VGND),
    .A1(_0867_),
    .A2(_1489_));
 sg13g2_nor2_2 _3568_ (.A(net842),
    .B(net847),
    .Y(_1490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3569_ (.B(_0877_),
    .C(_1490_),
    .A(_1972_),
    .Y(_1491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3570_ (.Y(_1492_),
    .A(net594),
    .B(_1491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3571_ (.A(net847),
    .B(net921),
    .C(net584),
    .Y(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3572_ (.Y(_1494_),
    .A(_0497_),
    .B(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3573_ (.Y(_0323_),
    .B1(net580),
    .B2(_1494_),
    .A2(net584),
    .A1(_1962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3574_ (.Y(_0324_),
    .B1(net580),
    .B2(_0497_),
    .A2(net584),
    .A1(_1963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3575_ (.Y(_1495_),
    .A(_0492_),
    .B(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3576_ (.Y(_0325_),
    .B1(net579),
    .B2(_1495_),
    .A2(_1492_),
    .A1(_1965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3577_ (.Y(_0326_),
    .B1(net579),
    .B2(_0494_),
    .A2(net583),
    .A1(_1964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3578_ (.Y(_0327_),
    .B1(net579),
    .B2(_0505_),
    .A2(net583),
    .A1(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3579_ (.Y(_0328_),
    .B1(net579),
    .B2(_0489_),
    .A2(net583),
    .A1(_1966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3580_ (.Y(_0329_),
    .B1(net579),
    .B2(_0496_),
    .A2(_1492_),
    .A1(_1969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3581_ (.Y(_0330_),
    .B1(net579),
    .B2(_0500_),
    .A2(net583),
    .A1(_1968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3582_ (.Y(_0331_),
    .B1(net580),
    .B2(_0498_),
    .A2(net584),
    .A1(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3583_ (.Y(_0332_),
    .B1(net580),
    .B2(_0499_),
    .A2(net584),
    .A1(_1959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3584_ (.Y(_0333_),
    .B1(net580),
    .B2(_1965_),
    .A2(net583),
    .A1(_1958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3585_ (.Y(_0334_),
    .B1(net579),
    .B2(_1964_),
    .A2(net583),
    .A1(_1957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3586_ (.Y(_0335_),
    .B1(_1493_),
    .B2(_1967_),
    .A2(net583),
    .A1(_1956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3587_ (.Y(_0336_),
    .B1(net580),
    .B2(_1966_),
    .A2(net584),
    .A1(_1955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3588_ (.Y(_0337_),
    .B1(net579),
    .B2(_1969_),
    .A2(net583),
    .A1(_1954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3589_ (.Y(_1496_),
    .A(_1968_),
    .B(_1494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3590_ (.Y(_0338_),
    .B1(net580),
    .B2(_1496_),
    .A2(net584),
    .A1(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3591_ (.Y(_1497_),
    .A(net488),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3592_ (.Y(_1498_),
    .B(_0549_),
    .A_N(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _3593_ (.A(net849),
    .B(_0551_),
    .C(_0552_),
    .Y(_1499_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_1498_));
 sg13g2_nor2b_2 _3594_ (.A(net777),
    .B_N(net774),
    .Y(_1500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3595_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net784),
    .A2(_0675_),
    .Y(_1501_),
    .B1(net783));
 sg13g2_nor2_1 _3596_ (.A(_0652_),
    .B(_1501_),
    .Y(_1502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3597_ (.Y(_1503_),
    .B(_1441_),
    .A_N(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3598_ (.Y(_1504_),
    .B(_1503_),
    .A_N(_0544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3599_ (.B1(_1500_),
    .VDD(VPWR),
    .Y(_1505_),
    .VSS(VGND),
    .A1(_1502_),
    .A2(_1504_));
 sg13g2_nand2_2 _3600_ (.Y(_1506_),
    .A(net780),
    .B(_0539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3601_ (.Y(_1507_),
    .A(_0539_),
    .B(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3602_ (.Y(_1508_),
    .B(_1507_),
    .A_N(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1506_),
    .A2(_1508_),
    .Y(_1509_),
    .B1(_0537_));
 sg13g2_nand2b_1 _3604_ (.Y(_1510_),
    .B(_0541_),
    .A_N(_0655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3605_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0647_),
    .A2(_0669_),
    .Y(_1511_),
    .B1(_1452_));
 sg13g2_nor2b_1 _3606_ (.A(net772),
    .B_N(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .Y(_1512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3607_ (.Y(_1513_),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .A_N(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3608_ (.A(net788),
    .B(net779),
    .C(_0539_),
    .Y(_1514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3609_ (.A(_0535_),
    .B(_0674_),
    .Y(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3610_ (.B1(_0545_),
    .VDD(VPWR),
    .Y(_1516_),
    .VSS(VGND),
    .A1(_1514_),
    .A2(_1515_));
 sg13g2_a21oi_1 _3611_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1510_),
    .A2(_1511_),
    .Y(_1517_),
    .B1(_1509_));
 sg13g2_nand4_1 _3612_ (.B(_1512_),
    .C(_1516_),
    .A(_1505_),
    .Y(_1518_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1517_));
 sg13g2_a22oi_1 _3613_ (.Y(_1519_),
    .B1(_1514_),
    .B2(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .A2(\u_usb_cdc.configured_o ),
    .A1(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3614_ (.A(net776),
    .B(_1926_),
    .Y(_1520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3615_ (.B(_0761_),
    .C(_1503_),
    .A(net783),
    .Y(_1521_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1520_));
 sg13g2_nand3_1 _3616_ (.B(_1519_),
    .C(_1521_),
    .A(_1518_),
    .Y(_1522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3617_ (.A(net753),
    .B(_1490_),
    .Y(_1523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3618_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1524_),
    .B(_1490_),
    .A(net753));
 sg13g2_nand2_1 _3619_ (.Y(_1525_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3620_ (.S0(net810),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .S1(net801),
    .X(_1526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3621_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net810),
    .A2(_1988_),
    .Y(_1527_),
    .B1(net801));
 sg13g2_o21ai_1 _3622_ (.B1(_1527_),
    .VDD(VPWR),
    .Y(_1528_),
    .VSS(VGND),
    .A1(net810),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ));
 sg13g2_mux2_1 _3623_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .S(net807),
    .X(_1529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3624_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_1529_),
    .Y(_1530_),
    .B1(_1923_));
 sg13g2_nand2_1 _3625_ (.Y(_1531_),
    .A(_1528_),
    .B(_1530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3626_ (.B1(_1531_),
    .VDD(VPWR),
    .Y(_1532_),
    .VSS(VGND),
    .A1(net797),
    .A2(_1526_));
 sg13g2_o21ai_1 _3627_ (.B1(_1525_),
    .VDD(VPWR),
    .Y(_1533_),
    .VSS(VGND),
    .A1(net795),
    .A2(_1532_));
 sg13g2_a221oi_1 _3628_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net637),
    .C1(net627),
    .B1(_1533_),
    .A1(_1499_),
    .Y(_1534_),
    .A2(_1522_));
 sg13g2_o21ai_1 _3629_ (.B1(net602),
    .VDD(VPWR),
    .Y(_1535_),
    .VSS(VGND),
    .A1(net187),
    .A2(_1523_));
 sg13g2_o21ai_1 _3630_ (.B1(_1497_),
    .VDD(VPWR),
    .Y(_0339_),
    .VSS(VGND),
    .A1(_1534_),
    .A2(_1535_));
 sg13g2_nand2_1 _3631_ (.Y(_1536_),
    .A(net560),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3632_ (.A(net784),
    .B(_0669_),
    .X(_1537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3633_ (.A(_0685_),
    .B(_1537_),
    .Y(_1538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3634_ (.A(_1538_),
    .B_N(net780),
    .Y(_1539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3635_ (.B(_1538_),
    .A(net780),
    .X(_1540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3636_ (.B(_0762_),
    .C(_1540_),
    .A(_0656_),
    .Y(_1541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3637_ (.Y(_1542_),
    .B(_1541_),
    .A_N(net773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3638_ (.B1(net781),
    .VDD(VPWR),
    .Y(_1543_),
    .VSS(VGND),
    .A1(net785),
    .A2(_1441_));
 sg13g2_o21ai_1 _3639_ (.B1(_0652_),
    .VDD(VPWR),
    .Y(_1544_),
    .VSS(VGND),
    .A1(net792),
    .A2(_0533_));
 sg13g2_o21ai_1 _3640_ (.B1(_1543_),
    .VDD(VPWR),
    .Y(_1545_),
    .VSS(VGND),
    .A1(net781),
    .A2(_1544_));
 sg13g2_a21oi_1 _3641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0533_),
    .A2(_1501_),
    .Y(_1546_),
    .B1(_1452_));
 sg13g2_o21ai_1 _3642_ (.B1(_1546_),
    .VDD(VPWR),
    .Y(_1547_),
    .VSS(VGND),
    .A1(_1441_),
    .A2(_1506_));
 sg13g2_a21oi_1 _3643_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1500_),
    .A2(_1545_),
    .Y(_1548_),
    .B1(_1513_));
 sg13g2_nand3_1 _3644_ (.B(_1547_),
    .C(_1548_),
    .A(_1542_),
    .Y(_1549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3645_ (.A(net779),
    .B(_0542_),
    .C(_0668_),
    .Y(_1550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3646_ (.Y(_1551_),
    .A(_1506_),
    .B(_1520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3647_ (.B1(_1549_),
    .VDD(VPWR),
    .Y(_1552_),
    .VSS(VGND),
    .A1(_1550_),
    .A2(_1551_));
 sg13g2_nand2_1 _3648_ (.Y(_1553_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3649_ (.S0(net806),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .S1(net799),
    .X(_1554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3650_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net807),
    .A2(_1989_),
    .Y(_1555_),
    .B1(net799));
 sg13g2_o21ai_1 _3651_ (.B1(_1555_),
    .VDD(VPWR),
    .Y(_1556_),
    .VSS(VGND),
    .A1(net807),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ));
 sg13g2_mux2_1 _3652_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .S(net807),
    .X(_1557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3653_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_1557_),
    .Y(_1558_),
    .B1(_1923_));
 sg13g2_nand2_1 _3654_ (.Y(_1559_),
    .A(_1556_),
    .B(_1558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3655_ (.B1(_1559_),
    .VDD(VPWR),
    .Y(_1560_),
    .VSS(VGND),
    .A1(net796),
    .A2(_1554_));
 sg13g2_o21ai_1 _3656_ (.B1(_1553_),
    .VDD(VPWR),
    .Y(_1561_),
    .VSS(VGND),
    .A1(net795),
    .A2(_1560_));
 sg13g2_a221oi_1 _3657_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net637),
    .C1(net627),
    .B1(_1561_),
    .A1(_1499_),
    .Y(_1562_),
    .A2(_1552_));
 sg13g2_o21ai_1 _3658_ (.B1(net602),
    .VDD(VPWR),
    .Y(_1563_),
    .VSS(VGND),
    .A1(net284),
    .A2(_1523_));
 sg13g2_o21ai_1 _3659_ (.B1(_1536_),
    .VDD(VPWR),
    .Y(_0340_),
    .VSS(VGND),
    .A1(_1562_),
    .A2(_1563_));
 sg13g2_a21o_1 _3660_ (.A2(_0762_),
    .A1(net781),
    .B1(_0544_),
    .X(_1564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3661_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0533_),
    .A2(_0541_),
    .Y(_1565_),
    .B1(net780));
 sg13g2_nor2_1 _3662_ (.A(net788),
    .B(_1506_),
    .Y(_1566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3663_ (.B1(net777),
    .VDD(VPWR),
    .Y(_1567_),
    .VSS(VGND),
    .A1(_1565_),
    .A2(_1566_));
 sg13g2_nor3_1 _3664_ (.A(net792),
    .B(_0533_),
    .C(_0657_),
    .Y(_1568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3665_ (.A(net773),
    .B(_1568_),
    .Y(_1569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3666_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net776),
    .A2(_0670_),
    .Y(_1570_),
    .B1(_0647_));
 sg13g2_a21oi_1 _3667_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0647_),
    .A2(_1441_),
    .Y(_1571_),
    .B1(_1570_));
 sg13g2_a21o_1 _3668_ (.A2(_1571_),
    .A1(net773),
    .B1(_1513_),
    .X(_1572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3669_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1569_),
    .C1(_1572_),
    .B1(_1567_),
    .A1(_1500_),
    .Y(_1573_),
    .A2(_1564_));
 sg13g2_nand2_1 _3670_ (.Y(_1574_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3671_ (.S0(net803),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .S1(net799),
    .X(_1575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3672_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net807),
    .A2(_1990_),
    .Y(_1576_),
    .B1(net799));
 sg13g2_o21ai_1 _3673_ (.B1(_1576_),
    .VDD(VPWR),
    .Y(_1577_),
    .VSS(VGND),
    .A1(net807),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ));
 sg13g2_mux2_1 _3674_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .S(net807),
    .X(_1578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3675_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_1578_),
    .Y(_1579_),
    .B1(_1923_));
 sg13g2_nand2_1 _3676_ (.Y(_1580_),
    .A(_1577_),
    .B(_1579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3677_ (.B1(_1580_),
    .VDD(VPWR),
    .Y(_1581_),
    .VSS(VGND),
    .A1(net796),
    .A2(_1575_));
 sg13g2_o21ai_1 _3678_ (.B1(_1574_),
    .VDD(VPWR),
    .Y(_1582_),
    .VSS(VGND),
    .A1(net795),
    .A2(_1581_));
 sg13g2_a221oi_1 _3679_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net637),
    .C1(net627),
    .B1(_1582_),
    .A1(_1499_),
    .Y(_1583_),
    .A2(_1573_));
 sg13g2_o21ai_1 _3680_ (.B1(net602),
    .VDD(VPWR),
    .Y(_1584_),
    .VSS(VGND),
    .A1(net232),
    .A2(_1523_));
 sg13g2_nand2_1 _3681_ (.Y(_1585_),
    .A(net519),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3682_ (.B1(_1585_),
    .VDD(VPWR),
    .Y(_0341_),
    .VSS(VGND),
    .A1(_1583_),
    .A2(_1584_));
 sg13g2_nand2_1 _3683_ (.Y(_1586_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3684_ (.A(net803),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .Y(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3685_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net803),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .Y(_1588_),
    .B1(_1587_));
 sg13g2_mux2_1 _3686_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .S(net803),
    .X(_1589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3687_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net799),
    .A2(_1589_),
    .Y(_1590_),
    .B1(net796));
 sg13g2_o21ai_1 _3688_ (.B1(_1590_),
    .VDD(VPWR),
    .Y(_1591_),
    .VSS(VGND),
    .A1(net799),
    .A2(_1588_));
 sg13g2_nor2b_1 _3689_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ),
    .B_N(net803),
    .Y(_1592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3690_ (.A(net803),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ),
    .Y(_1593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3691_ (.A(net799),
    .B(_1592_),
    .C(_1593_),
    .Y(_1594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3692_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .B_N(net803),
    .Y(_1595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3693_ (.B1(net799),
    .VDD(VPWR),
    .Y(_1596_),
    .VSS(VGND),
    .A1(net803),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ));
 sg13g2_o21ai_1 _3694_ (.B1(net796),
    .VDD(VPWR),
    .Y(_1597_),
    .VSS(VGND),
    .A1(_1595_),
    .A2(_1596_));
 sg13g2_o21ai_1 _3695_ (.B1(_1591_),
    .VDD(VPWR),
    .Y(_1598_),
    .VSS(VGND),
    .A1(_1594_),
    .A2(_1597_));
 sg13g2_o21ai_1 _3696_ (.B1(_1586_),
    .VDD(VPWR),
    .Y(_1599_),
    .VSS(VGND),
    .A1(net795),
    .A2(_1598_));
 sg13g2_nand3_1 _3697_ (.B(_1520_),
    .C(_1543_),
    .A(_0653_),
    .Y(_1600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3698_ (.A(net777),
    .B(_0658_),
    .Y(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3699_ (.Y(_1602_),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .B(_0537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3700_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .A2(_1507_),
    .Y(_1603_),
    .B1(_1602_));
 sg13g2_o21ai_1 _3701_ (.B1(_1603_),
    .VDD(VPWR),
    .Y(_1604_),
    .VSS(VGND),
    .A1(_0718_),
    .A2(_1601_));
 sg13g2_o21ai_1 _3702_ (.B1(net782),
    .VDD(VPWR),
    .Y(_1605_),
    .VSS(VGND),
    .A1(net792),
    .A2(net785));
 sg13g2_o21ai_1 _3703_ (.B1(_1500_),
    .VDD(VPWR),
    .Y(_1606_),
    .VSS(VGND),
    .A1(_1537_),
    .A2(_1605_));
 sg13g2_or2_1 _3704_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1607_),
    .B(_0685_),
    .A(net780));
 sg13g2_o21ai_1 _3705_ (.B1(_1606_),
    .VDD(VPWR),
    .Y(_1608_),
    .VSS(VGND),
    .A1(net773),
    .A2(_1607_));
 sg13g2_o21ai_1 _3706_ (.B1(_1600_),
    .VDD(VPWR),
    .Y(_1609_),
    .VSS(VGND),
    .A1(_1604_),
    .A2(_1608_));
 sg13g2_a221oi_1 _3707_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1499_),
    .C1(net627),
    .B1(_1609_),
    .A1(net637),
    .Y(_1610_),
    .A2(_1599_));
 sg13g2_o21ai_1 _3708_ (.B1(net602),
    .VDD(VPWR),
    .Y(_1611_),
    .VSS(VGND),
    .A1(net266),
    .A2(_1523_));
 sg13g2_nand2_1 _3709_ (.Y(_1612_),
    .A(net1005),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3710_ (.B1(_1612_),
    .VDD(VPWR),
    .Y(_0342_),
    .VSS(VGND),
    .A1(_1610_),
    .A2(_1611_));
 sg13g2_nand2_1 _3711_ (.Y(_1613_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3712_ (.A(net804),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .Y(_1614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3713_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net804),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .Y(_1615_),
    .B1(_1614_));
 sg13g2_mux2_1 _3714_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .S(net804),
    .X(_1616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3715_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net798),
    .A2(_1616_),
    .Y(_1617_),
    .B1(net796));
 sg13g2_o21ai_1 _3716_ (.B1(_1617_),
    .VDD(VPWR),
    .Y(_1618_),
    .VSS(VGND),
    .A1(net798),
    .A2(_1615_));
 sg13g2_nor2b_1 _3717_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ),
    .B_N(net805),
    .Y(_1619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3718_ (.A(net804),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ),
    .Y(_1620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3719_ (.A(net798),
    .B(_1619_),
    .C(_1620_),
    .Y(_1621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3720_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .B_N(net805),
    .Y(_1622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3721_ (.B1(net798),
    .VDD(VPWR),
    .Y(_1623_),
    .VSS(VGND),
    .A1(net805),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ));
 sg13g2_o21ai_1 _3722_ (.B1(net796),
    .VDD(VPWR),
    .Y(_1624_),
    .VSS(VGND),
    .A1(_1622_),
    .A2(_1623_));
 sg13g2_o21ai_1 _3723_ (.B1(_1618_),
    .VDD(VPWR),
    .Y(_1625_),
    .VSS(VGND),
    .A1(_1621_),
    .A2(_1624_));
 sg13g2_o21ai_1 _3724_ (.B1(_1613_),
    .VDD(VPWR),
    .Y(_1626_),
    .VSS(VGND),
    .A1(net795),
    .A2(_1625_));
 sg13g2_a21oi_1 _3725_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0545_),
    .A2(_0821_),
    .Y(_1627_),
    .B1(_1513_));
 sg13g2_o21ai_1 _3726_ (.B1(net773),
    .VDD(VPWR),
    .Y(_1628_),
    .VSS(VGND),
    .A1(_0543_),
    .A2(_0657_));
 sg13g2_a21oi_1 _3727_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0647_),
    .A2(_0674_),
    .Y(_1629_),
    .B1(_0537_));
 sg13g2_nand2_1 _3728_ (.Y(_1630_),
    .A(_1512_),
    .B(_1628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3729_ (.B(_1627_),
    .C(_1628_),
    .Y(_1631_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1629_));
 sg13g2_nand2_1 _3730_ (.Y(_1632_),
    .A(_1520_),
    .B(_1607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3731_ (.B1(_1631_),
    .VDD(VPWR),
    .Y(_1633_),
    .VSS(VGND),
    .A1(_1539_),
    .A2(_1632_));
 sg13g2_a221oi_1 _3732_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1499_),
    .C1(net627),
    .B1(_1633_),
    .A1(net637),
    .Y(_1634_),
    .A2(_1626_));
 sg13g2_o21ai_1 _3733_ (.B1(net602),
    .VDD(VPWR),
    .Y(_1635_),
    .VSS(VGND),
    .A1(net228),
    .A2(_1523_));
 sg13g2_nand2_1 _3734_ (.Y(_1636_),
    .A(net997),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3735_ (.B1(_1636_),
    .VDD(VPWR),
    .Y(_0343_),
    .VSS(VGND),
    .A1(_1634_),
    .A2(_1635_));
 sg13g2_nand2_1 _3736_ (.Y(_1637_),
    .A(net989),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3737_ (.Y(_1638_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3738_ (.A(net804),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .Y(_1639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3739_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net804),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .Y(_1640_),
    .B1(_1639_));
 sg13g2_mux2_1 _3740_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .S(net804),
    .X(_1641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3741_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net798),
    .A2(_1641_),
    .Y(_1642_),
    .B1(net796));
 sg13g2_o21ai_1 _3742_ (.B1(_1642_),
    .VDD(VPWR),
    .Y(_1643_),
    .VSS(VGND),
    .A1(net798),
    .A2(_1640_));
 sg13g2_nor2b_1 _3743_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ),
    .B_N(net805),
    .Y(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3744_ (.A(net808),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ),
    .Y(_1645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3745_ (.A(net798),
    .B(_1644_),
    .C(_1645_),
    .Y(_1646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3746_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .B_N(net805),
    .Y(_1647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3747_ (.B1(net800),
    .VDD(VPWR),
    .Y(_1648_),
    .VSS(VGND),
    .A1(net805),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ));
 sg13g2_o21ai_1 _3748_ (.B1(net796),
    .VDD(VPWR),
    .Y(_1649_),
    .VSS(VGND),
    .A1(_1647_),
    .A2(_1648_));
 sg13g2_o21ai_1 _3749_ (.B1(_1643_),
    .VDD(VPWR),
    .Y(_1650_),
    .VSS(VGND),
    .A1(_1646_),
    .A2(_1649_));
 sg13g2_o21ai_1 _3750_ (.B1(_1638_),
    .VDD(VPWR),
    .Y(_1651_),
    .VSS(VGND),
    .A1(net795),
    .A2(_1650_));
 sg13g2_or3_1 _3751_ (.A(_1926_),
    .B(_0533_),
    .C(_0657_),
    .X(_1652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3752_ (.Y(_1653_),
    .A(net866),
    .B(_1568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _3753_ (.A(net780),
    .B(_0543_),
    .C(_0761_),
    .D(_1503_),
    .X(_1654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3754_ (.A(net773),
    .B(_0544_),
    .C(_1654_),
    .Y(_1655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3755_ (.A(net776),
    .B_N(_1514_),
    .Y(_1656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3756_ (.B1(_1627_),
    .VDD(VPWR),
    .Y(_1657_),
    .VSS(VGND),
    .A1(_1628_),
    .A2(_1656_));
 sg13g2_o21ai_1 _3757_ (.B1(_1653_),
    .VDD(VPWR),
    .Y(_1658_),
    .VSS(VGND),
    .A1(_1655_),
    .A2(_1657_));
 sg13g2_a221oi_1 _3758_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1499_),
    .C1(net627),
    .B1(_1658_),
    .A1(net637),
    .Y(_1659_),
    .A2(_1651_));
 sg13g2_o21ai_1 _3759_ (.B1(net602),
    .VDD(VPWR),
    .Y(_1660_),
    .VSS(VGND),
    .A1(net236),
    .A2(_1523_));
 sg13g2_o21ai_1 _3760_ (.B1(_1637_),
    .VDD(VPWR),
    .Y(_0344_),
    .VSS(VGND),
    .A1(_1659_),
    .A2(_1660_));
 sg13g2_nand2_1 _3761_ (.Y(_1661_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .B(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _3762_ (.S0(net804),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .S1(net798),
    .X(_1662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3763_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net808),
    .A2(_1991_),
    .Y(_1663_),
    .B1(net800));
 sg13g2_o21ai_1 _3764_ (.B1(_1663_),
    .VDD(VPWR),
    .Y(_1664_),
    .VSS(VGND),
    .A1(net807),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ));
 sg13g2_mux2_1 _3765_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .S(net808),
    .X(_1665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3766_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_1665_),
    .Y(_1666_),
    .B1(_1923_));
 sg13g2_nand2_1 _3767_ (.Y(_1667_),
    .A(_1664_),
    .B(_1666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3768_ (.B1(_1667_),
    .VDD(VPWR),
    .Y(_1668_),
    .VSS(VGND),
    .A1(net797),
    .A2(_1662_));
 sg13g2_o21ai_1 _3769_ (.B1(_1661_),
    .VDD(VPWR),
    .Y(_1669_),
    .VSS(VGND),
    .A1(net795),
    .A2(_1668_));
 sg13g2_o21ai_1 _3770_ (.B1(_0537_),
    .VDD(VPWR),
    .Y(_1670_),
    .VSS(VGND),
    .A1(net773),
    .A2(_0536_));
 sg13g2_o21ai_1 _3771_ (.B1(_1652_),
    .VDD(VPWR),
    .Y(_1671_),
    .VSS(VGND),
    .A1(_1630_),
    .A2(_1670_));
 sg13g2_a221oi_1 _3772_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1499_),
    .C1(net627),
    .B1(_1671_),
    .A1(net638),
    .Y(_1672_),
    .A2(_1669_));
 sg13g2_o21ai_1 _3773_ (.B1(_0439_),
    .VDD(VPWR),
    .Y(_1673_),
    .VSS(VGND),
    .A1(net506),
    .A2(_1523_));
 sg13g2_nand2_1 _3774_ (.Y(_1674_),
    .A(net992),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3775_ (.B1(_1674_),
    .VDD(VPWR),
    .Y(_0345_),
    .VSS(VGND),
    .A1(_1672_),
    .A2(_1673_));
 sg13g2_a21oi_1 _3776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net810),
    .A2(_1992_),
    .Y(_1675_),
    .B1(net801));
 sg13g2_o21ai_1 _3777_ (.B1(_1675_),
    .VDD(VPWR),
    .Y(_1676_),
    .VSS(VGND),
    .A1(net810),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ));
 sg13g2_mux2_1 _3778_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .S(net808),
    .X(_1677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3779_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net801),
    .A2(_1677_),
    .Y(_1678_),
    .B1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ));
 sg13g2_nor2b_1 _3780_ (.A(net810),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .Y(_1679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3781_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net810),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .Y(_1680_),
    .B1(_1679_));
 sg13g2_mux2_1 _3782_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[63] ),
    .S(net808),
    .X(_1681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3783_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_1681_),
    .Y(_1682_),
    .B1(_1923_));
 sg13g2_o21ai_1 _3784_ (.B1(_1682_),
    .VDD(VPWR),
    .Y(_1683_),
    .VSS(VGND),
    .A1(net800),
    .A2(_1680_));
 sg13g2_a21oi_1 _3785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1676_),
    .A2(_1678_),
    .Y(_1684_),
    .B1(net795));
 sg13g2_a22oi_1 _3786_ (.Y(_1685_),
    .B1(_1683_),
    .B2(_1684_),
    .A2(net628),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[71] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3787_ (.VDD(VPWR),
    .Y(_1686_),
    .A(_1685_),
    .VSS(VGND));
 sg13g2_a22oi_1 _3788_ (.Y(_1687_),
    .B1(_1568_),
    .B2(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .A2(_1512_),
    .A1(_0660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3789_ (.VDD(VPWR),
    .Y(_1688_),
    .A(_1687_),
    .VSS(VGND));
 sg13g2_a221oi_1 _3790_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1499_),
    .C1(net627),
    .B1(_1688_),
    .A1(net637),
    .Y(_1689_),
    .A2(_1686_));
 sg13g2_o21ai_1 _3791_ (.B1(_0439_),
    .VDD(VPWR),
    .Y(_1690_),
    .VSS(VGND),
    .A1(net270),
    .A2(_1523_));
 sg13g2_nand2_1 _3792_ (.Y(_1691_),
    .A(net984),
    .B(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3793_ (.B1(_1691_),
    .VDD(VPWR),
    .Y(_0346_),
    .VSS(VGND),
    .A1(_1689_),
    .A2(_1690_));
 sg13g2_nand2_2 _3794_ (.Y(_1692_),
    .A(_1974_),
    .B(_0877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3795_ (.B(net592),
    .C(_1692_),
    .A(net767),
    .Y(_1693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3796_ (.B1(_1693_),
    .VDD(VPWR),
    .Y(_0347_),
    .VSS(VGND),
    .A1(net724),
    .A2(net600));
 sg13g2_nand3_1 _3797_ (.B(net592),
    .C(_1692_),
    .A(net766),
    .Y(_1694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3798_ (.B1(_1694_),
    .VDD(VPWR),
    .Y(_0348_),
    .VSS(VGND),
    .A1(net721),
    .A2(net600));
 sg13g2_nand3_1 _3799_ (.B(net592),
    .C(_1692_),
    .A(net765),
    .Y(_1695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3800_ (.B1(_1695_),
    .VDD(VPWR),
    .Y(_0349_),
    .VSS(VGND),
    .A1(_1913_),
    .A2(net600));
 sg13g2_nand3_1 _3801_ (.B(net592),
    .C(_1692_),
    .A(net1005),
    .Y(_1696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3802_ (.B1(_1696_),
    .VDD(VPWR),
    .Y(_0350_),
    .VSS(VGND),
    .A1(_1912_),
    .A2(net600));
 sg13g2_nand3_1 _3803_ (.B(net592),
    .C(_1692_),
    .A(net997),
    .Y(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3804_ (.B1(_1697_),
    .VDD(VPWR),
    .Y(_0351_),
    .VSS(VGND),
    .A1(_1915_),
    .A2(net600));
 sg13g2_nand3_1 _3805_ (.B(net592),
    .C(_1692_),
    .A(net989),
    .Y(_1698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3806_ (.B1(_1698_),
    .VDD(VPWR),
    .Y(_0352_),
    .VSS(VGND),
    .A1(_1914_),
    .A2(net600));
 sg13g2_nand3_1 _3807_ (.B(net592),
    .C(_1692_),
    .A(net992),
    .Y(_1699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3808_ (.B1(_1699_),
    .VDD(VPWR),
    .Y(_0353_),
    .VSS(VGND),
    .A1(_1917_),
    .A2(net600));
 sg13g2_nand3_1 _3809_ (.B(net592),
    .C(_1692_),
    .A(net984),
    .Y(_1700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3810_ (.B1(_1700_),
    .VDD(VPWR),
    .Y(_0354_),
    .VSS(VGND),
    .A1(_1916_),
    .A2(net600));
 sg13g2_nor2_2 _3811_ (.A(net841),
    .B(net847),
    .Y(_1701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3812_ (.Y(_1702_),
    .B1(_1701_),
    .B2(_1972_),
    .A2(_2017_),
    .A1(net848),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3813_ (.B(net593),
    .C(_0600_),
    .A(_0512_),
    .Y(_1703_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1702_));
 sg13g2_a21oi_1 _3814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_usb_cdc.ctrl_stall ),
    .A2(net641),
    .Y(_1704_),
    .B1(_0568_));
 sg13g2_nand2_1 _3815_ (.Y(_1705_),
    .A(net848),
    .B(_1704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3816_ (.B(_0862_),
    .C(_1701_),
    .A(net488),
    .Y(_1706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3817_ (.Y(_1707_),
    .A(_1705_),
    .B(_1706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3818_ (.A0(_1707_),
    .A1(net911),
    .S(_1703_),
    .X(_0355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3819_ (.Y(_1708_),
    .A(_0973_),
    .B(_1701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3820_ (.A0(_1708_),
    .A1(net944),
    .S(_1703_),
    .X(_0356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3821_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1709_),
    .B(_1701_),
    .A(_0517_));
 sg13g2_and2_1 _3822_ (.A(_0862_),
    .B(_1701_),
    .X(_1710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net765),
    .A2(_1710_),
    .Y(_1711_),
    .B1(_1703_));
 sg13g2_a22oi_1 _3824_ (.Y(_0357_),
    .B1(_1709_),
    .B2(_1711_),
    .A2(_1703_),
    .A1(_1934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3825_ (.A(_0990_),
    .B_N(_1704_),
    .Y(_1712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3826_ (.Y(_1713_),
    .B(net848),
    .A_N(_1712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3827_ (.Y(_1714_),
    .B1(net638),
    .B2(net771),
    .A2(net640),
    .A1(\u_usb_cdc.ctrl_stall ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3828_ (.VDD(VPWR),
    .Y(_1715_),
    .A(_1714_),
    .VSS(VGND));
 sg13g2_a221oi_1 _3829_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net841),
    .C1(_1703_),
    .B1(_1715_),
    .A1(net1005),
    .Y(_1716_),
    .A2(_1710_));
 sg13g2_a22oi_1 _3830_ (.Y(_0358_),
    .B1(_1713_),
    .B2(_1716_),
    .A2(_1703_),
    .A1(_1935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3831_ (.A0(_0436_),
    .A1(_0603_),
    .S(_1474_),
    .X(_1717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3832_ (.A(net717),
    .B(_1717_),
    .Y(_1718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3833_ (.VDD(VPWR),
    .Y(_1719_),
    .A(_1718_),
    .VSS(VGND));
 sg13g2_nor3_1 _3834_ (.A(net840),
    .B(_0436_),
    .C(_1474_),
    .Y(_1720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3835_ (.B1(net756),
    .VDD(VPWR),
    .Y(_1721_),
    .VSS(VGND),
    .A1(_1719_),
    .A2(_1720_));
 sg13g2_nor2_1 _3836_ (.A(_0510_),
    .B(_0956_),
    .Y(_1722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3837_ (.B1(_0713_),
    .VDD(VPWR),
    .Y(_1723_),
    .VSS(VGND),
    .A1(_0506_),
    .A2(_1722_));
 sg13g2_nand4_1 _3838_ (.B(net745),
    .C(_0437_),
    .A(net840),
    .Y(_1724_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1723_));
 sg13g2_nand2_1 _3839_ (.Y(_0359_),
    .A(_1721_),
    .B(_1724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3840_ (.A(net752),
    .B(net717),
    .C(_0436_),
    .D(_0950_),
    .Y(_1725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _3841_ (.A(_1934_),
    .B(_0450_),
    .C(_0452_),
    .D(_0481_),
    .X(_1726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3842_ (.B1(_1726_),
    .VDD(VPWR),
    .Y(_1727_),
    .VSS(VGND),
    .A1(_0578_),
    .A2(_0956_));
 sg13g2_a21oi_1 _3843_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1725_),
    .A2(_1727_),
    .Y(_1728_),
    .B1(net107));
 sg13g2_a21oi_1 _3844_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1474_),
    .A2(_1718_),
    .Y(_0360_),
    .B1(_1728_));
 sg13g2_o21ai_1 _3845_ (.B1(_0912_),
    .VDD(VPWR),
    .Y(_1729_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .A2(_0905_));
 sg13g2_nand3_1 _3846_ (.B(_0899_),
    .C(_1729_),
    .A(net312),
    .Y(_1730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3847_ (.B1(_1730_),
    .VDD(VPWR),
    .Y(_0361_),
    .VSS(VGND),
    .A1(_1946_),
    .A2(net595));
 sg13g2_nand3_1 _3848_ (.B(_0899_),
    .C(_1729_),
    .A(net209),
    .Y(_1731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3849_ (.B1(_1731_),
    .VDD(VPWR),
    .Y(_0362_),
    .VSS(VGND),
    .A1(_1947_),
    .A2(net595));
 sg13g2_nand3_1 _3850_ (.B(_0899_),
    .C(_1729_),
    .A(net421),
    .Y(_1732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3851_ (.B1(_1732_),
    .VDD(VPWR),
    .Y(_0363_),
    .VSS(VGND),
    .A1(_1949_),
    .A2(net595));
 sg13g2_nand3_1 _3852_ (.B(_0899_),
    .C(_1729_),
    .A(net329),
    .Y(_1733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3853_ (.B1(_1733_),
    .VDD(VPWR),
    .Y(_0364_),
    .VSS(VGND),
    .A1(_1948_),
    .A2(net595));
 sg13g2_nand3_1 _3854_ (.B(_0899_),
    .C(_1729_),
    .A(net310),
    .Y(_1734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3855_ (.B1(_1734_),
    .VDD(VPWR),
    .Y(_0365_),
    .VSS(VGND),
    .A1(_1951_),
    .A2(net595));
 sg13g2_nand3_1 _3856_ (.B(_0899_),
    .C(_1729_),
    .A(net338),
    .Y(_1735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3857_ (.B1(_1735_),
    .VDD(VPWR),
    .Y(_0366_),
    .VSS(VGND),
    .A1(_1950_),
    .A2(net595));
 sg13g2_nand3_1 _3858_ (.B(_0899_),
    .C(_1729_),
    .A(net496),
    .Y(_1736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3859_ (.B1(_1736_),
    .VDD(VPWR),
    .Y(_0367_),
    .VSS(VGND),
    .A1(_1952_),
    .A2(net595));
 sg13g2_nand2_1 _3860_ (.Y(_1737_),
    .A(_0056_),
    .B(_1946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3861_ (.B(_0884_),
    .C(_1737_),
    .A(_0883_),
    .Y(_1738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3862_ (.A2(_1738_),
    .A1(_0889_),
    .B1(_0906_),
    .X(_1739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3863_ (.B(\u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .C(net961),
    .Y(_1740_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0056_));
 sg13g2_o21ai_1 _3864_ (.B1(_1739_),
    .VDD(VPWR),
    .Y(_1741_),
    .VSS(VGND),
    .A1(_2039_),
    .A2(net962));
 sg13g2_mux2_1 _3865_ (.A0(net496),
    .A1(net963),
    .S(_0901_),
    .X(_0368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3866_ (.A(_0901_),
    .B_N(net1039),
    .Y(_1742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3867_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net1007),
    .C1(_2039_),
    .B1(_0898_),
    .A1(_2044_),
    .Y(_1743_),
    .A2(_0881_));
 sg13g2_or2_1 _3868_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0369_),
    .B(_1743_),
    .A(_1742_));
 sg13g2_nor2_2 _3869_ (.A(_1978_),
    .B(_2003_),
    .Y(_1744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3870_ (.A(\u_usb_cdc.u_sie.u_phy_rx.state_q[1] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ),
    .C(_1744_),
    .Y(_1745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3871_ (.A(net713),
    .B(_1745_),
    .Y(_1746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3872_ (.Y(_1747_),
    .B(net744),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1745_));
 sg13g2_nor2_1 _3873_ (.A(net361),
    .B(net615),
    .Y(_1748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3874_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net741),
    .A2(net361),
    .Y(_0370_),
    .B1(_1748_));
 sg13g2_a21oi_1 _3875_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net361),
    .A2(net365),
    .Y(_1749_),
    .B1(_1745_));
 sg13g2_nor2_1 _3876_ (.A(net716),
    .B(_1749_),
    .Y(_1750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3877_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net741),
    .A2(net361),
    .Y(_1751_),
    .B1(net365));
 sg13g2_nor2_1 _3878_ (.A(_1750_),
    .B(net366),
    .Y(_0371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3879_ (.B1(net336),
    .VDD(VPWR),
    .Y(_1752_),
    .VSS(VGND),
    .A1(net716),
    .A2(_1749_));
 sg13g2_nand3_1 _3880_ (.B(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .C(net615),
    .A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .Y(_1753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3881_ (.B1(_1752_),
    .VDD(VPWR),
    .Y(_0372_),
    .VSS(VGND),
    .A1(net336),
    .A2(_1753_));
 sg13g2_and4_1 _3882_ (.A(net361),
    .B(net365),
    .C(net336),
    .D(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .X(_1754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3883_ (.B1(net741),
    .VDD(VPWR),
    .Y(_1755_),
    .VSS(VGND),
    .A1(_1745_),
    .A2(_1754_));
 sg13g2_nand4_1 _3884_ (.B(net361),
    .C(net365),
    .A(net741),
    .Y(_1756_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net336));
 sg13g2_nand2b_1 _3885_ (.Y(_1757_),
    .B(_1756_),
    .A_N(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3886_ (.A(_1755_),
    .B(_1757_),
    .X(_0373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3887_ (.Y(_1758_),
    .A(net348),
    .B(_1755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3888_ (.Y(_1759_),
    .A(net615),
    .B(_1754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3889_ (.B1(_1758_),
    .VDD(VPWR),
    .Y(_0374_),
    .VSS(VGND),
    .A1(net348),
    .A2(_1759_));
 sg13g2_and3_2 _3890_ (.X(_1760_),
    .A(net348),
    .B(net387),
    .C(_1754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3891_ (.A(_1745_),
    .B(_1760_),
    .Y(_1761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3892_ (.A(net713),
    .B(_1761_),
    .Y(_1762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3893_ (.B(net348),
    .C(_1754_),
    .A(net741),
    .Y(_1763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3894_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2004_),
    .A2(_1763_),
    .Y(_0375_),
    .B1(_1762_));
 sg13g2_a21oi_1 _3895_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net615),
    .A2(_1760_),
    .Y(_1764_),
    .B1(net282));
 sg13g2_a21oi_1 _3896_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net282),
    .A2(_1762_),
    .Y(_0376_),
    .B1(_1764_));
 sg13g2_and3_1 _3897_ (.X(_1765_),
    .A(net282),
    .B(net879),
    .C(_1760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3898_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net282),
    .A2(_1760_),
    .Y(_1766_),
    .B1(net879));
 sg13g2_nor3_1 _3899_ (.A(_1747_),
    .B(_1765_),
    .C(_1766_),
    .Y(_1767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3900_ (.A2(net879),
    .A1(net713),
    .B1(_1767_),
    .X(_0377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3901_ (.Y(_1768_),
    .A(net713),
    .B(net457),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3902_ (.A(net457),
    .B(_1765_),
    .X(_1769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3903_ (.B1(net615),
    .VDD(VPWR),
    .Y(_1770_),
    .VSS(VGND),
    .A1(net457),
    .A2(_1765_));
 sg13g2_o21ai_1 _3904_ (.B1(_1768_),
    .VDD(VPWR),
    .Y(_0378_),
    .VSS(VGND),
    .A1(_1769_),
    .A2(_1770_));
 sg13g2_nand2_1 _3905_ (.Y(_1771_),
    .A(net714),
    .B(net391),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3906_ (.A(net391),
    .B(_1769_),
    .X(_1772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3907_ (.B1(net615),
    .VDD(VPWR),
    .Y(_1773_),
    .VSS(VGND),
    .A1(net391),
    .A2(_1769_));
 sg13g2_o21ai_1 _3908_ (.B1(_1771_),
    .VDD(VPWR),
    .Y(_0379_),
    .VSS(VGND),
    .A1(_1772_),
    .A2(_1773_));
 sg13g2_nand2_1 _3909_ (.Y(_1774_),
    .A(net714),
    .B(net340),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3910_ (.A(net340),
    .B(_1772_),
    .X(_1775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3911_ (.B1(net615),
    .VDD(VPWR),
    .Y(_1776_),
    .VSS(VGND),
    .A1(net340),
    .A2(_1772_));
 sg13g2_o21ai_1 _3912_ (.B1(_1774_),
    .VDD(VPWR),
    .Y(_0380_),
    .VSS(VGND),
    .A1(_1775_),
    .A2(_1776_));
 sg13g2_nand2_1 _3913_ (.Y(_1777_),
    .A(net713),
    .B(net437),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3914_ (.Y(_1778_),
    .A(net437),
    .B(_1775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3915_ (.B1(_1777_),
    .VDD(VPWR),
    .Y(_0381_),
    .VSS(VGND),
    .A1(_1747_),
    .A2(_1778_));
 sg13g2_a21oi_1 _3916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net437),
    .A2(_1775_),
    .Y(_1779_),
    .B1(net896));
 sg13g2_and3_1 _3917_ (.X(_1780_),
    .A(net437),
    .B(net896),
    .C(_1775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3918_ (.A(_1747_),
    .B(_1779_),
    .C(_1780_),
    .Y(_1781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3919_ (.A2(net896),
    .A1(net713),
    .B1(_1781_),
    .X(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3920_ (.Y(_1782_),
    .A(net713),
    .B(net319),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3921_ (.A(net319),
    .B(_1780_),
    .X(_1783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3922_ (.B1(net615),
    .VDD(VPWR),
    .Y(_1784_),
    .VSS(VGND),
    .A1(net319),
    .A2(_1780_));
 sg13g2_o21ai_1 _3923_ (.B1(_1782_),
    .VDD(VPWR),
    .Y(_0383_),
    .VSS(VGND),
    .A1(_1783_),
    .A2(_1784_));
 sg13g2_nand2_1 _3924_ (.Y(_1785_),
    .A(net714),
    .B(net352),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3925_ (.A(net352),
    .B(_1783_),
    .X(_1786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3926_ (.B1(_1746_),
    .VDD(VPWR),
    .Y(_1787_),
    .VSS(VGND),
    .A1(net352),
    .A2(_1783_));
 sg13g2_o21ai_1 _3927_ (.B1(_1785_),
    .VDD(VPWR),
    .Y(_0384_),
    .VSS(VGND),
    .A1(_1786_),
    .A2(_1787_));
 sg13g2_nand2_1 _3928_ (.Y(_1788_),
    .A(net714),
    .B(net353),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3929_ (.A(net353),
    .B(_1786_),
    .X(_1789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3930_ (.B1(_1746_),
    .VDD(VPWR),
    .Y(_1790_),
    .VSS(VGND),
    .A1(net353),
    .A2(_1786_));
 sg13g2_o21ai_1 _3931_ (.B1(_1788_),
    .VDD(VPWR),
    .Y(_0385_),
    .VSS(VGND),
    .A1(_1789_),
    .A2(_1790_));
 sg13g2_nand2_1 _3932_ (.Y(_1791_),
    .A(net717),
    .B(net853),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3933_ (.A(net853),
    .B(_1789_),
    .Y(_1792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3934_ (.A2(_1789_),
    .A1(net853),
    .B1(_1747_),
    .X(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3935_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1791_),
    .A2(_1793_),
    .Y(_0386_),
    .B1(_1792_));
 sg13g2_nand3_1 _3936_ (.B(_1746_),
    .C(_1789_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .Y(_1794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3937_ (.Y(_0387_),
    .B1(_1794_),
    .B2(_1976_),
    .A2(_1793_),
    .A1(_0916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3938_ (.Y(_1795_),
    .A(_2037_),
    .B(_0904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3939_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0910_),
    .A2(_1795_),
    .Y(_1796_),
    .B1(_0909_));
 sg13g2_mux2_1 _3940_ (.A0(_1796_),
    .A1(net707),
    .S(net979),
    .X(_0388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3941_ (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .X(_1797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3942_ (.Y(_1798_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .B(net423),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3943_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1796_),
    .A2(_1798_),
    .Y(_1799_),
    .B1(net707));
 sg13g2_a21oi_1 _3944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .A2(_1796_),
    .Y(_1800_),
    .B1(net423));
 sg13g2_nor2_1 _3945_ (.A(_1799_),
    .B(net424),
    .Y(_0389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3946_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1796_),
    .A2(_1797_),
    .Y(_1801_),
    .B1(net57));
 sg13g2_a21oi_1 _3947_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net57),
    .A2(_1799_),
    .Y(_0390_),
    .B1(_1801_));
 sg13g2_nor2_1 _3948_ (.A(net713),
    .B(_1744_),
    .Y(_1802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3949_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net744),
    .A2(net387),
    .Y(_1803_),
    .B1(net917));
 sg13g2_nor2_1 _3950_ (.A(_1802_),
    .B(net918),
    .Y(_0391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3951_ (.A(net465),
    .B(net747),
    .Y(_1804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3952_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net747),
    .A2(_0945_),
    .Y(_0392_),
    .B1(_1804_));
 sg13g2_nor2_1 _3953_ (.A(net754),
    .B(net747),
    .Y(_1805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3954_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net747),
    .A2(net306),
    .Y(_0393_),
    .B1(_1805_));
 sg13g2_nor2_2 _3955_ (.A(net955),
    .B(net413),
    .Y(_1806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3956_ (.A(_1978_),
    .B(net368),
    .C(net708),
    .D(_1806_),
    .Y(_1807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3957_ (.A2(net708),
    .A1(net976),
    .B1(_1807_),
    .X(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3958_ (.A(net751),
    .B(net746),
    .Y(_1808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3959_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net746),
    .A2(_0943_),
    .Y(_0395_),
    .B1(_1808_));
 sg13g2_nor2_1 _3960_ (.A(net553),
    .B(_2040_),
    .Y(_1809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3961_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1943_),
    .A2(_2040_),
    .Y(_0396_),
    .B1(net554));
 sg13g2_nor2_1 _3962_ (.A(net556),
    .B(_2040_),
    .Y(_1810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3963_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1944_),
    .A2(_2040_),
    .Y(_0397_),
    .B1(net557));
 sg13g2_nor2_1 _3964_ (.A(net452),
    .B(net708),
    .Y(_1811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3965_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1943_),
    .A2(net708),
    .Y(_0398_),
    .B1(net453));
 sg13g2_nor2_1 _3966_ (.A(net532),
    .B(net708),
    .Y(_1812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3967_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1944_),
    .A2(net708),
    .Y(_0399_),
    .B1(net533));
 sg13g2_o21ai_1 _3968_ (.B1(_0988_),
    .VDD(VPWR),
    .Y(_0400_),
    .VSS(VGND),
    .A1(_1918_),
    .A2(net742));
 sg13g2_nand2_1 _3969_ (.Y(_1813_),
    .A(net187),
    .B(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3970_ (.B1(_1813_),
    .VDD(VPWR),
    .Y(_0401_),
    .VSS(VGND),
    .A1(_1947_),
    .A2(net614));
 sg13g2_nand2_1 _3971_ (.Y(_1814_),
    .A(net284),
    .B(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3972_ (.B1(net285),
    .VDD(VPWR),
    .Y(_0402_),
    .VSS(VGND),
    .A1(_1949_),
    .A2(net614));
 sg13g2_nand2_1 _3973_ (.Y(_1815_),
    .A(net232),
    .B(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3974_ (.B1(_1815_),
    .VDD(VPWR),
    .Y(_0403_),
    .VSS(VGND),
    .A1(_1948_),
    .A2(net613));
 sg13g2_nand2_1 _3975_ (.Y(_1816_),
    .A(net266),
    .B(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3976_ (.B1(_1816_),
    .VDD(VPWR),
    .Y(_0404_),
    .VSS(VGND),
    .A1(_1951_),
    .A2(net613));
 sg13g2_nand2_1 _3977_ (.Y(_1817_),
    .A(net228),
    .B(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3978_ (.B1(_1817_),
    .VDD(VPWR),
    .Y(_0405_),
    .VSS(VGND),
    .A1(_1950_),
    .A2(net613));
 sg13g2_nand2_1 _3979_ (.Y(_1818_),
    .A(net236),
    .B(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3980_ (.B1(_1818_),
    .VDD(VPWR),
    .Y(_0406_),
    .VSS(VGND),
    .A1(_1952_),
    .A2(net613));
 sg13g2_mux2_1 _3981_ (.A0(net496),
    .A1(net506),
    .S(net614),
    .X(_0407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3982_ (.Y(_1819_),
    .A(net270),
    .B(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3983_ (.B1(_1819_),
    .VDD(VPWR),
    .Y(_0408_),
    .VSS(VGND),
    .A1(_0056_),
    .A2(net614));
 sg13g2_nor2_1 _3984_ (.A(net748),
    .B(net885),
    .Y(_1820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3985_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net748),
    .A2(_0921_),
    .Y(_0409_),
    .B1(net886));
 sg13g2_a22oi_1 _3986_ (.Y(_1821_),
    .B1(_0433_),
    .B2(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .A2(_2027_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3987_ (.B1(_1821_),
    .VDD(VPWR),
    .Y(_1822_),
    .VSS(VGND),
    .A1(_1921_),
    .A2(net709));
 sg13g2_nor2_2 _3988_ (.A(net754),
    .B(_0925_),
    .Y(_1823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3989_ (.Y(_1824_),
    .B1(net767),
    .B2(net842),
    .A2(\u_usb_cdc.u_sie.pid_q[0] ),
    .A1(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3990_ (.Y(_1825_),
    .B1(_1968_),
    .B2(net837),
    .A2(_1953_),
    .A1(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3991_ (.B(_1824_),
    .C(_1825_),
    .A(_1705_),
    .Y(_1826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3992_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1823_),
    .A2(_1826_),
    .Y(_1827_),
    .B1(_1822_));
 sg13g2_nor2_1 _3993_ (.A(net904),
    .B(net709),
    .Y(_1828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3994_ (.A(_1008_),
    .B(_1827_),
    .C(_1828_),
    .X(_1829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3995_ (.A(_2020_),
    .B(_1008_),
    .X(_1830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3996_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net904),
    .A2(_1830_),
    .Y(_1831_),
    .B1(net643));
 sg13g2_a22oi_1 _3997_ (.Y(_0410_),
    .B1(_1829_),
    .B2(_1831_),
    .A2(net643),
    .A1(_1993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3998_ (.A(_2027_),
    .B(_0925_),
    .Y(_1832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3999_ (.Y(_1833_),
    .A(net709),
    .B(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4000_ (.B1(net709),
    .VDD(VPWR),
    .Y(_1834_),
    .VSS(VGND),
    .A1(net835),
    .A2(_0926_));
 sg13g2_nor2_1 _4001_ (.A(_2027_),
    .B(_1008_),
    .Y(_1835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4002_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1836_),
    .VSS(VGND),
    .A1(net439),
    .A2(_1835_));
 sg13g2_a22oi_1 _4003_ (.Y(_1837_),
    .B1(_1969_),
    .B2(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .A2(net766),
    .A1(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4004_ (.Y(_1838_),
    .B1(_1954_),
    .B2(net845),
    .A2(\u_usb_cdc.u_sie.pid_q[1] ),
    .A1(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4005_ (.B(_1837_),
    .C(_1838_),
    .A(_2018_),
    .Y(_1839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0926_),
    .A2(_1839_),
    .Y(_1840_),
    .B1(_1834_));
 sg13g2_nor4_1 _4007_ (.A(_2028_),
    .B(_1009_),
    .C(_1836_),
    .D(_1840_),
    .Y(_1841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4008_ (.A2(net642),
    .A1(net904),
    .B1(_1841_),
    .X(_0411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4009_ (.A(net642),
    .B(_1009_),
    .Y(_1842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4010_ (.Y(_1843_),
    .B1(_1955_),
    .B2(net845),
    .A2(\u_usb_cdc.u_sie.pid_q[2] ),
    .A1(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4011_ (.Y(_1844_),
    .B1(_1966_),
    .B2(net837),
    .A2(net765),
    .A1(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4012_ (.B(_1843_),
    .C(_1844_),
    .A(_0518_),
    .Y(_1845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4013_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0926_),
    .A2(_1845_),
    .Y(_1846_),
    .B1(_1834_));
 sg13g2_o21ai_1 _4014_ (.B1(_1842_),
    .VDD(VPWR),
    .Y(_1847_),
    .VSS(VGND),
    .A1(net383),
    .A2(_1835_));
 sg13g2_nor3_1 _4015_ (.A(_2028_),
    .B(_1846_),
    .C(_1847_),
    .Y(_1848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4016_ (.A2(net642),
    .A1(net439),
    .B1(_1848_),
    .X(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4017_ (.Y(_1849_),
    .B1(_1956_),
    .B2(net845),
    .A2(\u_usb_cdc.u_sie.pid_q[3] ),
    .A1(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4018_ (.Y(_1850_),
    .B1(_1967_),
    .B2(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .A2(\u_usb_cdc.u_sie.data_q[3] ),
    .A1(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4019_ (.A(net626),
    .B(_2026_),
    .C(_1849_),
    .D(_1850_),
    .X(_1851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4020_ (.B1(_1851_),
    .VDD(VPWR),
    .Y(_1852_),
    .VSS(VGND),
    .A1(_2018_),
    .A2(_1712_));
 sg13g2_nand2_1 _4021_ (.Y(_1853_),
    .A(_1979_),
    .B(_2028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4022_ (.Y(_1854_),
    .B(_2027_),
    .A_N(net292),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4023_ (.B(_1852_),
    .C(_1853_),
    .A(_0926_),
    .Y(_1855_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1854_));
 sg13g2_a21o_1 _4024_ (.A2(_2027_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .B1(_1830_),
    .X(_1856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4025_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net292),
    .A2(_1856_),
    .Y(_1857_),
    .B1(net642));
 sg13g2_a22oi_1 _4026_ (.Y(_0413_),
    .B1(_1855_),
    .B2(_1857_),
    .A2(net642),
    .A1(_1994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4027_ (.Y(_1858_),
    .A(net292),
    .B(net643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4028_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1859_),
    .B(_1704_),
    .A(_2018_));
 sg13g2_a22oi_1 _4029_ (.Y(_1860_),
    .B1(_1957_),
    .B2(net845),
    .A2(_1932_),
    .A1(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4030_ (.Y(_1861_),
    .B1(_1964_),
    .B2(net837),
    .A2(\u_usb_cdc.u_sie.data_q[4] ),
    .A1(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4031_ (.B(_1860_),
    .C(_1861_),
    .A(_1859_),
    .Y(_1862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4032_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1823_),
    .C1(_1822_),
    .B1(_1862_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .Y(_1863_),
    .A2(_1830_));
 sg13g2_o21ai_1 _4033_ (.B1(net625),
    .VDD(VPWR),
    .Y(_1864_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .A2(_2026_));
 sg13g2_o21ai_1 _4034_ (.B1(_1858_),
    .VDD(VPWR),
    .Y(_0414_),
    .VSS(VGND),
    .A1(_1863_),
    .A2(_1864_));
 sg13g2_nand2_1 _4035_ (.Y(_1865_),
    .A(net356),
    .B(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4036_ (.Y(_1866_),
    .B1(_1965_),
    .B2(net837),
    .A2(_1958_),
    .A1(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4037_ (.Y(_1867_),
    .B1(\u_usb_cdc.u_sie.data_q[5] ),
    .B2(net843),
    .A2(_1933_),
    .A1(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4038_ (.Y(_1868_),
    .A(_1866_),
    .B(_1867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4039_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1868_),
    .C1(_1834_),
    .B1(_1823_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .Y(_1869_),
    .A2(_0433_));
 sg13g2_o21ai_1 _4040_ (.B1(_1842_),
    .VDD(VPWR),
    .Y(_1870_),
    .VSS(VGND),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .A2(_1835_));
 sg13g2_o21ai_1 _4041_ (.B1(_1865_),
    .VDD(VPWR),
    .Y(_0415_),
    .VSS(VGND),
    .A1(_1869_),
    .A2(_1870_));
 sg13g2_a22oi_1 _4042_ (.Y(_1871_),
    .B1(_1963_),
    .B2(net837),
    .A2(_1934_),
    .A1(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4043_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net842),
    .C1(_0570_),
    .B1(\u_usb_cdc.u_sie.data_q[6] ),
    .A1(net845),
    .Y(_1872_),
    .A2(_1959_));
 sg13g2_nand2_1 _4044_ (.Y(_1873_),
    .A(_1871_),
    .B(_1872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4045_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1823_),
    .A2(_1873_),
    .Y(_1874_),
    .B1(_1834_));
 sg13g2_a22oi_1 _4046_ (.Y(_1875_),
    .B1(_1874_),
    .B2(_1821_),
    .A2(_1834_),
    .A1(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4047_ (.Y(_1876_),
    .B1(_1842_),
    .B2(_1875_),
    .A2(net642),
    .A1(net494),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4048_ (.VDD(VPWR),
    .Y(_0416_),
    .A(net495),
    .VSS(VGND));
 sg13g2_nand2_1 _4049_ (.Y(_1877_),
    .A(net848),
    .B(_1712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4050_ (.Y(_1878_),
    .B1(_1961_),
    .B2(net845),
    .A2(_1935_),
    .A1(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4051_ (.Y(_1879_),
    .B1(_1962_),
    .B2(net837),
    .A2(\u_usb_cdc.u_sie.data_q[7] ),
    .A1(net843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4052_ (.B(_1877_),
    .C(_1878_),
    .A(net626),
    .Y(_1880_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1879_));
 sg13g2_a22oi_1 _4053_ (.Y(_1881_),
    .B1(_1832_),
    .B2(_1880_),
    .A2(net709),
    .A1(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4054_ (.Y(_1882_),
    .B1(_1842_),
    .B2(_1881_),
    .A2(net642),
    .A1(net459),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4055_ (.VDD(VPWR),
    .Y(_0417_),
    .A(net460),
    .VSS(VGND));
 sg13g2_nor2_1 _4056_ (.A(net308),
    .B(_1842_),
    .Y(_1883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4057_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net308),
    .A2(_2023_),
    .Y(_0418_),
    .B1(_1883_));
 sg13g2_nor2_1 _4058_ (.A(net643),
    .B(_1010_),
    .Y(_1884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4059_ (.B(_0922_),
    .A(net937),
    .X(_1885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4060_ (.A(_1884_),
    .B(_1885_),
    .Y(_0419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4061_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0059_),
    .A2(net308),
    .Y(_1886_),
    .B1(net481));
 sg13g2_nor2_1 _4062_ (.A(_1884_),
    .B(_1886_),
    .Y(_1887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _4063_ (.A(net835),
    .B(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .C(_2020_),
    .D(_1833_),
    .Y(_1888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4064_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0923_),
    .A2(_1887_),
    .Y(_1889_),
    .B1(_1888_));
 sg13g2_a21oi_1 _4065_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1908_),
    .A2(net643),
    .Y(_0420_),
    .B1(_1889_));
 sg13g2_nand3_1 _4066_ (.B(_2036_),
    .C(_0882_),
    .A(net748),
    .Y(_1890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4067_ (.B1(_1890_),
    .VDD(VPWR),
    .Y(_0421_),
    .VSS(VGND),
    .A1(net748),
    .A2(_2003_));
 sg13g2_nand2_1 _4068_ (.Y(_1891_),
    .A(_1979_),
    .B(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4069_ (.B(net625),
    .C(_1853_),
    .A(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .Y(_1892_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1891_));
 sg13g2_nand2_1 _4070_ (.Y(_1893_),
    .A(net350),
    .B(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4071_ (.B1(_1893_),
    .VDD(VPWR),
    .Y(_0422_),
    .VSS(VGND),
    .A1(net350),
    .A2(_1892_));
 sg13g2_nand2_1 _4072_ (.Y(_1894_),
    .A(net389),
    .B(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4073_ (.Y(_1895_),
    .A(net350),
    .B(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4074_ (.B1(_1894_),
    .VDD(VPWR),
    .Y(_0423_),
    .VSS(VGND),
    .A1(_1892_),
    .A2(_1895_));
 sg13g2_nand2_1 _4075_ (.Y(_1896_),
    .A(net404),
    .B(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4076_ (.Y(_1897_),
    .A(net350),
    .B(net389),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4077_ (.B(_1897_),
    .A(net404),
    .X(_1898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4078_ (.B1(_1896_),
    .VDD(VPWR),
    .Y(_0424_),
    .VSS(VGND),
    .A1(_1892_),
    .A2(_1898_));
 sg13g2_nor3_1 _4079_ (.A(net598),
    .B(_0586_),
    .C(_1524_),
    .Y(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4080_ (.Y(_1900_),
    .A(net638),
    .B(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4081_ (.Y(_1901_),
    .A(net84),
    .B(_1900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4082_ (.B1(_1901_),
    .VDD(VPWR),
    .Y(_0425_),
    .VSS(VGND),
    .A1(_1919_),
    .A2(_1900_));
 sg13g2_nand2_1 _4083_ (.Y(_1902_),
    .A(net640),
    .B(_1899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4084_ (.Y(_1903_),
    .A(net164),
    .B(_1902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4085_ (.B1(_1903_),
    .VDD(VPWR),
    .Y(_0426_),
    .VSS(VGND),
    .A1(_1919_),
    .A2(_1902_));
 sg13g2_mux2_1 _4086_ (.A0(_1023_),
    .A1(net834),
    .S(_1031_),
    .X(_1904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4087_ (.A0(net884),
    .A1(_1904_),
    .S(_1128_),
    .X(_0427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4088_ (.Y(_1905_),
    .A(net547),
    .B(_1031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4089_ (.B(net647),
    .C(_1905_),
    .A(net749),
    .Y(_1906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4090_ (.B1(_1906_),
    .VDD(VPWR),
    .Y(_1907_),
    .VSS(VGND),
    .A1(net749),
    .A2(net551));
 sg13g2_inv_1 _4091_ (.VDD(VPWR),
    .Y(_0428_),
    .A(net552),
    .VSS(VGND));
 sg13g2_buf_1 _4092_ (.A(_0053_),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _4093_ (.RESET_B(net689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net487),
    .Q(\u_usb_cdc.u_sie.out_toggle_q[0] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _4094_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net939),
    .Q(_0048_),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_2 _4095_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net895),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_2 _4096_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net867),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4097_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net943),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _4098_ (.RESET_B(net689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net875),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _4099_ (.RESET_B(net690),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net514),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _4100_ (.RESET_B(net689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net484),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_2 _4101_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net958),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_2 _4102_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net975),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4103_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0010_),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4104_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net412),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4105_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net523),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4106_ (.RESET_B(net689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net56),
    .Q(\u_usb_cdc.u_sie.out_toggle_q[1] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _4107_ (.RESET_B(net688),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net407),
    .Q(\u_usb_cdc.u_sie.in_toggle_q[0] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _4108_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net858),
    .Q(\u_usb_cdc.u_sie.in_toggle_q[1] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _4109_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net380),
    .Q(\u_usb_cdc.u_sie.in_toggle_q[2] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _4110_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net542),
    .Q(_0049_),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _4111_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net960),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _4112_ (.RESET_B(net689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0012_),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _4113_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net970),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _4114_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0014_),
    .Q(\u_usb_cdc.ctrl_stall ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _4115_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net472),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[5] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _4116_ (.RESET_B(net694),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net948),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _4117_ (.RESET_B(net694),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net950),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _4118_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0063_),
    .Q(_0050_),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _4119_ (.RESET_B(net699),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0020_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[1] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _4120_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net525),
    .Q(\u_usb_cdc.u_sie.phy_state_q[2] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4121_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0022_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[3] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4122_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0023_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[4] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _4123_ (.RESET_B(net688),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net302),
    .Q(\u_usb_cdc.u_sie.phy_state_q[5] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _4124_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net142),
    .Q(\u_usb_cdc.u_sie.phy_state_q[6] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _4125_ (.RESET_B(net698),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0026_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[7] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _4126_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0027_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[8] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4127_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net505),
    .Q(\u_usb_cdc.u_sie.phy_state_q[9] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _4128_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0018_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _4129_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0019_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _4130_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1023),
    .Q(_0051_),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _4131_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net574),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _4132_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1008),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _4133_ (.RESET_B(net736),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0031_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _4134_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net315),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _4135_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0065_),
    .Q(_0052_),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _4136_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net395),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.state_q[1] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _4137_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0034_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _4138_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net930),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.state_q[3] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _4139_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net263),
    .Q(\u_usb_cdc.u_sie.addr_q[0] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _4140_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0066_),
    .Q(_0053_),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _4141_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _4142_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net369),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _4143_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0038_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _4144_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net300),
    .Q(_0054_),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _4145_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net548),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _4146_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0075_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _4147_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0076_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _4148_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _4149_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _4150_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0079_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _4151_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _4152_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _4153_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _4154_ (.RESET_B(net680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net462),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4155_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net550),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _4156_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net491),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _4157_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net434),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _4158_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net444),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _4159_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net456),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _4160_ (.RESET_B(net664),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net527),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4161_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net870),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _4162_ (.RESET_B(net680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net83),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4163_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net194),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _4164_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net77),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _4165_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net79),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _4166_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net120),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _4167_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net132),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _4168_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net221),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4169_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net106),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _4170_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net251),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4171_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net169),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _4172_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net183),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _4173_ (.RESET_B(net665),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net249),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _4174_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net95),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _4175_ (.RESET_B(net664),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net73),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _4176_ (.RESET_B(net670),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net239),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4177_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net122),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4178_ (.RESET_B(net680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net516),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4179_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net512),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _4180_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net538),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _4181_ (.RESET_B(net665),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net529),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _4182_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net536),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _4183_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net521),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _4184_ (.RESET_B(net664),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net571),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _4185_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net510),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _4186_ (.RESET_B(net680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net159),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4187_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net219),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4188_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net155),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4189_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net199),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4190_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net206),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4191_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net114),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4192_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net197),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4193_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net178),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _4194_ (.RESET_B(net680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net63),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4195_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net65),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4196_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net75),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _4197_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net60),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _4198_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net91),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _4199_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net118),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4200_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net71),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4201_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net97),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _4202_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net89),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4203_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net81),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4204_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net254),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _4205_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net87),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _4206_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net136),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _4207_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net241),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4208_ (.RESET_B(net670),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net243),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4209_ (.RESET_B(net670),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net151),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4210_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net508),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4211_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net518),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4212_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net470),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4213_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net468),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4214_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net476),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4215_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net464),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4216_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net480),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _4217_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net478),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[63] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4218_ (.RESET_B(net680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net93),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4219_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net201),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4220_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net110),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _4221_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net124),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4222_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net134),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _4223_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net140),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4224_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net69),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _4225_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net138),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[71] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _4226_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net860),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _4227_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net863),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _4228_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net883),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _4229_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\u_usb_cdc.in_ready_o [0]),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _4230_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net978),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _4231_ (.RESET_B(net679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0160_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _4232_ (.RESET_B(net679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _4233_ (.RESET_B(net679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _4234_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _4235_ (.RESET_B(net679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net852),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _4236_ (.RESET_B(net679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net420),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _4237_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net364),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _4238_ (.RESET_B(net675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net217),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4239_ (.RESET_B(net675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4240_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net289),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4241_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[3] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4242_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4243_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net287),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4244_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net256),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[6] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4245_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0174_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4246_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net204),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4247_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net104),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4248_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net67),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4249_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net279),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[11] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4250_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net112),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4251_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net269),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4252_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net223),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[14] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4253_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net116),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _4254_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net399),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4255_ (.RESET_B(net655),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net442),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4256_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net326),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[18] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4257_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net332),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4258_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4259_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net360),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4260_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net346),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4261_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net335),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[23] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4262_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net173),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4263_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4264_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net291),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[26] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4265_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4266_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net281),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[28] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4267_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net273),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[29] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4268_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net161),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4269_ (.RESET_B(net674),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net371),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[31] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4270_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net258),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4271_ (.RESET_B(net655),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net144),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4272_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net181),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4273_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net126),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[35] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4274_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net186),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4275_ (.RESET_B(net655),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net190),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4276_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net247),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[38] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4277_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net213),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4278_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net215),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4279_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net147),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4280_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net176),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4281_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net128),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4282_ (.RESET_B(net655),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net231),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4283_ (.RESET_B(net655),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net163),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _4284_ (.RESET_B(net650),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net235),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4285_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net99),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4286_ (.RESET_B(net675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net318),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4287_ (.RESET_B(net675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net344),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4288_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net417),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4289_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0218_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[51] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4290_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0219_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4291_ (.RESET_B(net674),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net403),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4292_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net427),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[54] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4293_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4294_ (.RESET_B(net675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net225),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4295_ (.RESET_B(net675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net102),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4296_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net277),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4297_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[59] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4298_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4299_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net324),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4300_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net373),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[62] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4301_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net149),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4302_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net153),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[64] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4303_ (.RESET_B(net650),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net130),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[65] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4304_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net208),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[66] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4305_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net192),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[67] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4306_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0235_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[68] ),
    .CLK(clknet_3_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _4307_ (.RESET_B(net650),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net227),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[69] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4308_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net167),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[70] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4309_ (.RESET_B(net650),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net171),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[71] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4310_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0239_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _4311_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net893),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _4312_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0241_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _4313_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0242_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _4314_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0243_),
    .Q(net19),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4315_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net297),
    .Q(net20),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4316_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net260),
    .Q(net21),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4317_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net447),
    .Q(net22),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4318_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net52),
    .Q(net23),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4319_ (.RESET_B(net651),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net245),
    .Q(net24),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4320_ (.RESET_B(net651),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net295),
    .Q(net25),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _4321_ (.RESET_B(net651),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net265),
    .Q(net26),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4322_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1004),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _4323_ (.RESET_B(net653),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net936),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _4324_ (.RESET_B(net653),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net941),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _4325_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net952),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _4326_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net544),
    .Q(\u_usb_cdc.out_valid_o [0]),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _4327_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0255_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _4328_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[1] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _4329_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1032),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _4330_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net966),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4331_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0259_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[0] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _4332_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1016),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[1] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _4333_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0261_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _4334_ (.RESET_B(net682),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net981),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _4335_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0263_),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[0] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _4336_ (.RESET_B(net685),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[1] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _4337_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net546),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[2] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _4338_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0266_),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[3] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _4339_ (.RESET_B(net685),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0267_),
    .Q(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _4340_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0268_),
    .Q(\u_usb_cdc.addr[0] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _4341_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0269_),
    .Q(\u_usb_cdc.addr[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _4342_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0270_),
    .Q(\u_usb_cdc.addr[2] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _4343_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0271_),
    .Q(\u_usb_cdc.addr[3] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _4344_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0272_),
    .Q(\u_usb_cdc.addr[4] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _4345_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0273_),
    .Q(\u_usb_cdc.addr[5] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _4346_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0274_),
    .Q(\u_usb_cdc.addr[6] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4347_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0275_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[0] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4348_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0276_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[1] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4349_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net429),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[2] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4350_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0278_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[3] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4351_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0279_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[4] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4352_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net474),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[5] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4353_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net436),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[6] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4354_ (.RESET_B(net690),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0282_),
    .Q(_0055_),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _4355_ (.RESET_B(net690),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0283_),
    .Q(\u_usb_cdc.u_ctrl_endp.dev_state_q[1] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_2 _4356_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0284_),
    .Q(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _4357_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net954),
    .Q(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _4358_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net493),
    .Q(\u_usb_cdc.u_ctrl_endp.class_q ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _4359_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0287_),
    .Q(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4360_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0288_),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _4361_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net927),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4362_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net865),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4363_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net899),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _4364_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0292_),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _4365_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net909),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _4366_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net565),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _4367_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0295_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _4368_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0296_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _4369_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0297_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _4370_ (.RESET_B(net694),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0298_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _4371_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0299_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _4372_ (.RESET_B(net694),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0300_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _4373_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net563),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _4374_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0302_),
    .Q(\u_usb_cdc.bulk_out_nak [0]),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _4375_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0303_),
    .Q(\u_usb_cdc.endp[0] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _4376_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0304_),
    .Q(\u_usb_cdc.endp[1] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _4377_ (.RESET_B(net688),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0305_),
    .Q(\u_usb_cdc.endp[2] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _4378_ (.RESET_B(net688),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0306_),
    .Q(\u_usb_cdc.endp[3] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _4379_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0307_),
    .Q(\u_usb_cdc.u_sie.addr_q[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _4380_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net386),
    .Q(\u_usb_cdc.u_sie.addr_q[2] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4381_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0309_),
    .Q(\u_usb_cdc.u_sie.addr_q[3] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4382_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0310_),
    .Q(\u_usb_cdc.u_sie.addr_q[4] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4383_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net382),
    .Q(\u_usb_cdc.u_sie.addr_q[5] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _4384_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net410),
    .Q(\u_usb_cdc.u_sie.addr_q[6] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _4385_ (.RESET_B(net728),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net956),
    .Q(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_2 _4386_ (.RESET_B(net728),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net415),
    .Q(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_2 _4387_ (.RESET_B(net699),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0315_),
    .Q(\u_usb_cdc.sie_in_req ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _4388_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net355),
    .Q(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _4389_ (.RESET_B(net698),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net432),
    .Q(\u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _4390_ (.RESET_B(net698),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net157),
    .Q(\u_usb_cdc.u_sie.delay_cnt_q[2] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _4391_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net328),
    .Q(\u_usb_cdc.u_sie.in_byte_q[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _4392_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net377),
    .Q(\u_usb_cdc.u_sie.in_byte_q[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4393_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net322),
    .Q(\u_usb_cdc.u_sie.in_byte_q[2] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4394_ (.RESET_B(net698),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net401),
    .Q(\u_usb_cdc.u_sie.in_byte_q[3] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4395_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net531),
    .Q(\u_usb_cdc.u_sie.crc16_q[0] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4396_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0324_),
    .Q(\u_usb_cdc.u_sie.crc16_q[1] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4397_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0325_),
    .Q(\u_usb_cdc.u_sie.crc16_q[2] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4398_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0326_),
    .Q(\u_usb_cdc.u_sie.crc16_q[3] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4399_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0327_),
    .Q(\u_usb_cdc.u_sie.crc16_q[4] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4400_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0328_),
    .Q(\u_usb_cdc.u_sie.crc16_q[5] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4401_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net907),
    .Q(\u_usb_cdc.u_sie.crc16_q[6] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4402_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net891),
    .Q(\u_usb_cdc.u_sie.crc16_q[7] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4403_ (.RESET_B(net696),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net916),
    .Q(\u_usb_cdc.u_sie.crc16_q[8] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _4404_ (.RESET_B(net696),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net889),
    .Q(\u_usb_cdc.u_sie.crc16_q[9] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _4405_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net855),
    .Q(\u_usb_cdc.u_sie.crc16_q[10] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _4406_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net903),
    .Q(\u_usb_cdc.u_sie.crc16_q[11] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4407_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net914),
    .Q(\u_usb_cdc.u_sie.crc16_q[12] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _4408_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net540),
    .Q(\u_usb_cdc.u_sie.crc16_q[13] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4409_ (.RESET_B(net696),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0337_),
    .Q(\u_usb_cdc.u_sie.crc16_q[14] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4410_ (.RESET_B(net696),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0338_),
    .Q(\u_usb_cdc.u_sie.crc16_q[15] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _4411_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0339_),
    .Q(\u_usb_cdc.u_sie.data_q[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _4412_ (.RESET_B(net706),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0340_),
    .Q(\u_usb_cdc.u_sie.data_q[1] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _4413_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0341_),
    .Q(\u_usb_cdc.u_sie.data_q[2] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _4414_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0342_),
    .Q(\u_usb_cdc.u_sie.data_q[3] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _4415_ (.RESET_B(net694),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0343_),
    .Q(\u_usb_cdc.u_sie.data_q[4] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _4416_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0344_),
    .Q(\u_usb_cdc.u_sie.data_q[5] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _4417_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0345_),
    .Q(\u_usb_cdc.u_sie.data_q[6] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _4418_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0346_),
    .Q(\u_usb_cdc.u_sie.data_q[7] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4419_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0347_),
    .Q(\u_usb_cdc.sie_out_data[0] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _4420_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0348_),
    .Q(\u_usb_cdc.sie_out_data[1] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _4421_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0349_),
    .Q(\u_usb_cdc.sie_out_data[2] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _4422_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0350_),
    .Q(\u_usb_cdc.sie_out_data[3] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _4423_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0351_),
    .Q(\u_usb_cdc.sie_out_data[4] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _4424_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0352_),
    .Q(\u_usb_cdc.sie_out_data[5] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _4425_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0353_),
    .Q(\u_usb_cdc.sie_out_data[6] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _4426_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0354_),
    .Q(\u_usb_cdc.sie_out_data[7] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _4427_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net912),
    .Q(\u_usb_cdc.u_sie.pid_q[0] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _4428_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net945),
    .Q(\u_usb_cdc.u_sie.pid_q[1] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _4429_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net999),
    .Q(\u_usb_cdc.u_sie.pid_q[2] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _4430_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1029),
    .Q(\u_usb_cdc.u_sie.pid_q[3] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _4431_ (.RESET_B(net699),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0359_),
    .Q(\u_usb_cdc.sie_out_err ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _4432_ (.RESET_B(net699),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net108),
    .Q(\u_usb_cdc.u_sie.out_eop_q ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _4433_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net313),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _4434_ (.RESET_B(net731),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net210),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _4435_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net422),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[2] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _4436_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net330),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _4437_ (.RESET_B(net731),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net311),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _4438_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net339),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[5] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _4439_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net497),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _4440_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net964),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _4441_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0369_),
    .Q(_0056_),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _4442_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net362),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_2 _4443_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net367),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _4444_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net337),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _4445_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net983),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _4446_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net349),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4447_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net388),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _4448_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net283),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _4449_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0377_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4450_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net458),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _4451_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net392),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4452_ (.RESET_B(net726),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net341),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _4453_ (.RESET_B(net726),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net438),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4454_ (.RESET_B(net726),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0382_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4455_ (.RESET_B(net726),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net320),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4456_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0384_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4457_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0385_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _4458_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0386_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _4459_ (.RESET_B(net728),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net275),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _4460_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0388_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _4461_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net425),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _4462_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net58),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _4463_ (.RESET_B(net726),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net919),
    .Q(\u_usb_cdc.bus_reset ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _4464_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net466),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4465_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net877),
    .Q(\u_usb_cdc.u_sie.rx_err ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _4466_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0394_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _4467_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net503),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_q ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _4468_ (.RESET_B(net732),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0395_),
    .Q(\u_usb_cdc.u_sie.rx_valid ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4469_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net307),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_err_q ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _4470_ (.RESET_B(net736),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net555),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _4471_ (.RESET_B(net736),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net558),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _4472_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net454),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _4473_ (.RESET_B(net736),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net534),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _4474_ (.RESET_B(net689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0400_),
    .Q(\u_usb_cdc.sie_in_data_ack ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _4475_ (.RESET_B(net732),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net451),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_valid_q ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4476_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net188),
    .Q(\u_usb_cdc.u_sie.rx_data[0] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _4477_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0402_),
    .Q(\u_usb_cdc.u_sie.rx_data[1] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _4478_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net233),
    .Q(\u_usb_cdc.u_sie.rx_data[2] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _4479_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net267),
    .Q(\u_usb_cdc.u_sie.rx_data[3] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _4480_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net229),
    .Q(\u_usb_cdc.u_sie.rx_data[4] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _4481_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net237),
    .Q(\u_usb_cdc.u_sie.rx_data[5] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _4482_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0407_),
    .Q(\u_usb_cdc.u_sie.rx_data[6] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4483_ (.RESET_B(net732),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net271),
    .Q(\u_usb_cdc.u_sie.rx_data[7] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4484_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net54),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[0] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4485_ (.RESET_B(net737),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0047_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[1] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _4486_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net887),
    .Q(net31),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _4487_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net47),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4488_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net46),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _4489_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net13),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _4490_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net48),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4491_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net44),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4492_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net12),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _4493_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0410_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _4494_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0411_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _4495_ (.RESET_B(net701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0412_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[2] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _4496_ (.RESET_B(net701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net384),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[3] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _4497_ (.RESET_B(net701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net293),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _4498_ (.RESET_B(net701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net357),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _4499_ (.RESET_B(net701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0416_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _4500_ (.RESET_B(net701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0417_),
    .Q(_0057_),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _4501_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net309),
    .Q(_0058_),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _4502_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0419_),
    .Q(_0059_),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _4503_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net482),
    .Q(_0060_),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _4504_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net375),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.se0_q ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _4505_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net351),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _4506_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net390),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4507_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net405),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4508_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\u_usb_cdc.clk_gate_q ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _4509_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0039_),
    .Q(\u_usb_cdc.clk_cnt_q[0] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _4510_ (.RESET_B(net731),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0040_),
    .Q(\u_usb_cdc.clk_cnt_q[1] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _4511_ (.RESET_B(net1),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net45),
    .Q(\u_usb_cdc.rstn ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _4512_ (.RESET_B(net1),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net38),
    .Q(\u_usb_cdc.rstn_sq[1] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _4513_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net85),
    .Q(\u_usb_cdc.u_sie.in_zlp_q[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4514_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net165),
    .Q(\u_usb_cdc.u_sie.in_zlp_q[0] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4515_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0427_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _4516_ (.RESET_B(net679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0428_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_tiehi heichips25_usb_cdc_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi heichips25_usb_cdc_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi heichips25_usb_cdc_41 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi heichips25_usb_cdc_42 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi heichips25_usb_cdc_43 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_usb_cdc_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net33));
 sg13g2_tielo heichips25_usb_cdc_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net34));
 sg13g2_tielo heichips25_usb_cdc_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net35));
 sg13g2_tielo heichips25_usb_cdc_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net36));
 sg13g2_tielo heichips25_usb_cdc_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net37));
 sg13g2_tiehi _4512__38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_buf_1 _4529_ (.A(\u_usb_cdc.out_valid_o [0]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4530_ (.A(\u_usb_cdc.in_ready_o [0]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 _4531_ (.A(\u_usb_cdc.configured_o ),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _4532_ (.A(net27),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 spad_env_f_bit i_spad_env_f_bit (.VGND(VGND),
    .VPWR(VPWR),
    .clk(clknet_1_0__leaf_clk),
    .env_bit(net18),
    .env_valid(net14),
    .spad_hit_async(uio_in[2]));
 sg13g2_buf_2 fanout576 (.A(_1419_),
    .X(net576),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout577 (.A(_1419_),
    .X(net577),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout578 (.A(_1390_),
    .X(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout579 (.A(net580),
    .X(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout580 (.A(_1493_),
    .X(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout581 (.A(_1401_),
    .X(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout582 (.A(_1401_),
    .X(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout583 (.A(net584),
    .X(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout584 (.A(_1492_),
    .X(net584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout585 (.A(net587),
    .X(net585),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout586 (.A(net587),
    .X(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout587 (.A(_1002_),
    .X(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout588 (.A(_0622_),
    .X(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout589 (.A(_0622_),
    .X(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout590 (.A(_0618_),
    .X(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout591 (.A(_0618_),
    .X(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout592 (.A(net594),
    .X(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout593 (.A(net594),
    .X(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout594 (.A(_0521_),
    .X(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout595 (.A(_0901_),
    .X(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout596 (.A(net599),
    .X(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout597 (.A(net599),
    .X(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout598 (.A(net599),
    .X(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout599 (.A(_0440_),
    .X(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout600 (.A(net602),
    .X(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout601 (.A(net602),
    .X(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout602 (.A(_0439_),
    .X(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout603 (.A(net604),
    .X(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout604 (.A(_1232_),
    .X(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout605 (.A(net607),
    .X(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout606 (.A(net607),
    .X(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout607 (.A(_1195_),
    .X(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout608 (.A(net609),
    .X(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout609 (.A(_1204_),
    .X(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout610 (.A(net612),
    .X(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout611 (.A(net612),
    .X(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout612 (.A(_1099_),
    .X(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout613 (.A(net614),
    .X(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout614 (.A(_0942_),
    .X(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout615 (.A(_1746_),
    .X(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout617 (.A(_1284_),
    .X(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout618 (.A(net621),
    .X(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout619 (.A(net621),
    .X(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout620 (.A(net621),
    .X(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout621 (.A(_1044_),
    .X(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout622 (.A(net623),
    .X(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout623 (.A(_0697_),
    .X(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout624 (.A(_0630_),
    .X(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout625 (.A(_2023_),
    .X(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout626 (.A(_2020_),
    .X(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout627 (.A(_1524_),
    .X(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout628 (.A(_1371_),
    .X(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout629 (.A(_1294_),
    .X(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout630 (.A(net631),
    .X(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout631 (.A(_1222_),
    .X(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout632 (.A(net633),
    .X(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout633 (.A(_1176_),
    .X(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout634 (.A(net635),
    .X(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout635 (.A(_1142_),
    .X(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout636 (.A(_1078_),
    .X(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout637 (.A(net638),
    .X(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout639 (.A(_0567_),
    .X(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout640 (.A(net641),
    .X(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout641 (.A(_0515_),
    .X(net641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout642 (.A(net643),
    .X(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout643 (.A(_2024_),
    .X(net643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout644 (.A(_1059_),
    .X(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout645 (.A(_1039_),
    .X(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout646 (.A(net647),
    .X(net646),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout647 (.A(_1014_),
    .X(net647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout648 (.A(net651),
    .X(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout649 (.A(net651),
    .X(net649),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout651 (.A(net653),
    .X(net651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout652 (.A(net653),
    .X(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout653 (.A(net671),
    .X(net653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout654 (.A(net659),
    .X(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout655 (.A(net659),
    .X(net655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout656 (.A(net659),
    .X(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout657 (.A(net659),
    .X(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout658 (.A(net659),
    .X(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout659 (.A(net671),
    .X(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout660 (.A(net661),
    .X(net660),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout661 (.A(net665),
    .X(net661),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout662 (.A(net664),
    .X(net662),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout663 (.A(net665),
    .X(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout665 (.A(net671),
    .X(net665),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout666 (.A(net667),
    .X(net666),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout667 (.A(net671),
    .X(net667),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout668 (.A(net670),
    .X(net668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout669 (.A(net670),
    .X(net669),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout670 (.A(net671),
    .X(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout671 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ),
    .X(net671),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout672 (.A(net674),
    .X(net672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout673 (.A(net674),
    .X(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout674 (.A(net675),
    .X(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout675 (.A(net682),
    .X(net675),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout676 (.A(net682),
    .X(net676),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout677 (.A(net682),
    .X(net677),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout678 (.A(net680),
    .X(net678),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout679 (.A(net680),
    .X(net679),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout680 (.A(net682),
    .X(net680),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout681 (.A(net682),
    .X(net681),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout682 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ),
    .X(net682),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout683 (.A(net685),
    .X(net683),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout684 (.A(net685),
    .X(net684),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout685 (.A(net690),
    .X(net685),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout686 (.A(net690),
    .X(net686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout687 (.A(net689),
    .X(net687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout688 (.A(net689),
    .X(net688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout689 (.A(net690),
    .X(net689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout690 (.A(net706),
    .X(net690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout691 (.A(net692),
    .X(net691),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout692 (.A(net706),
    .X(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout693 (.A(net694),
    .X(net693),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout694 (.A(net706),
    .X(net694),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout695 (.A(net704),
    .X(net695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout696 (.A(net704),
    .X(net696),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout697 (.A(net699),
    .X(net697),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout698 (.A(net699),
    .X(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout699 (.A(net704),
    .X(net699),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout700 (.A(net704),
    .X(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout701 (.A(net704),
    .X(net701),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout703 (.A(net704),
    .X(net703),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout704 (.A(net705),
    .X(net704),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout705 (.A(net706),
    .X(net705),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout706 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ),
    .X(net706),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout707 (.A(net708),
    .X(net707),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout708 (.A(_2041_),
    .X(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout709 (.A(_2026_),
    .X(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout710 (.A(_2015_),
    .X(net710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout711 (.A(_1980_),
    .X(net711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout712 (.A(_1980_),
    .X(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout713 (.A(net715),
    .X(net713),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout714 (.A(net715),
    .X(net714),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout715 (.A(net716),
    .X(net715),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout716 (.A(_1939_),
    .X(net716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout717 (.A(_1939_),
    .X(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout718 (.A(_1939_),
    .X(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout719 (.A(_1916_),
    .X(net719),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout720 (.A(_1912_),
    .X(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout721 (.A(net722),
    .X(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout722 (.A(_1911_),
    .X(net722),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout723 (.A(_1910_),
    .X(net723),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout724 (.A(_1910_),
    .X(net724),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout725 (.A(net738),
    .X(net725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout726 (.A(net738),
    .X(net726),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout727 (.A(net728),
    .X(net727),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout728 (.A(net738),
    .X(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout729 (.A(net731),
    .X(net729),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout730 (.A(net731),
    .X(net730),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout731 (.A(net732),
    .X(net731),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout732 (.A(net738),
    .X(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout733 (.A(net734),
    .X(net733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout734 (.A(net737),
    .X(net734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout735 (.A(net737),
    .X(net735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout736 (.A(net737),
    .X(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout737 (.A(net738),
    .X(net737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout738 (.A(net1048),
    .X(net738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout739 (.A(net741),
    .X(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout740 (.A(net741),
    .X(net740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout741 (.A(net749),
    .X(net741),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout742 (.A(net743),
    .X(net742),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout743 (.A(net744),
    .X(net743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout744 (.A(net749),
    .X(net744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout745 (.A(net746),
    .X(net745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout746 (.A(net747),
    .X(net746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout747 (.A(net748),
    .X(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout748 (.A(net749),
    .X(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout749 (.A(\u_usb_cdc.clk_gate_q ),
    .X(net749),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout750 (.A(net751),
    .X(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout751 (.A(net934),
    .X(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout752 (.A(net753),
    .X(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout753 (.A(net754),
    .X(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout754 (.A(net876),
    .X(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout755 (.A(net1043),
    .X(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout756 (.A(net1043),
    .X(net756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout757 (.A(net1012),
    .X(net757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout758 (.A(net1024),
    .X(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout759 (.A(net298),
    .X(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout760 (.A(net1033),
    .X(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout761 (.A(net1045),
    .X(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout762 (.A(\u_usb_cdc.sie_out_data[1] ),
    .X(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout763 (.A(net764),
    .X(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout764 (.A(\u_usb_cdc.sie_out_data[0] ),
    .X(net764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout765 (.A(net519),
    .X(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout766 (.A(net560),
    .X(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout767 (.A(net488),
    .X(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout768 (.A(net769),
    .X(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout769 (.A(\u_usb_cdc.endp[0] ),
    .X(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout770 (.A(net771),
    .X(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout771 (.A(\u_usb_cdc.bulk_out_nak [0]),
    .X(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout772 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .X(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout773 (.A(net775),
    .X(net773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout774 (.A(net775),
    .X(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout775 (.A(net1049),
    .X(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout776 (.A(net778),
    .X(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout777 (.A(net778),
    .X(net777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout778 (.A(net1021),
    .X(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout779 (.A(net783),
    .X(net779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout780 (.A(net781),
    .X(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout781 (.A(net782),
    .X(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout782 (.A(net783),
    .X(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout783 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .X(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout784 (.A(net786),
    .X(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout785 (.A(net786),
    .X(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout786 (.A(net787),
    .X(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout787 (.A(net1050),
    .X(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout788 (.A(net789),
    .X(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout789 (.A(net790),
    .X(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout790 (.A(net1052),
    .X(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout791 (.A(net793),
    .X(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout792 (.A(net793),
    .X(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout793 (.A(net1011),
    .X(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout794 (.A(net946),
    .X(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout795 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .X(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout796 (.A(net797),
    .X(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout797 (.A(net1040),
    .X(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout798 (.A(net800),
    .X(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout799 (.A(net800),
    .X(net799),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout800 (.A(net802),
    .X(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout801 (.A(net802),
    .X(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout802 (.A(net1014),
    .X(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout803 (.A(net806),
    .X(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout804 (.A(net806),
    .X(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout805 (.A(net806),
    .X(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout806 (.A(net811),
    .X(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout807 (.A(net811),
    .X(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout808 (.A(net811),
    .X(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout809 (.A(net810),
    .X(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout810 (.A(net811),
    .X(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout811 (.A(net1038),
    .X(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout812 (.A(net813),
    .X(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout813 (.A(net1031),
    .X(net813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout814 (.A(net817),
    .X(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout815 (.A(net817),
    .X(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout816 (.A(net817),
    .X(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout817 (.A(net1051),
    .X(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout818 (.A(net819),
    .X(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout819 (.A(net820),
    .X(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout820 (.A(net1041),
    .X(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout821 (.A(net825),
    .X(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout822 (.A(net823),
    .X(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout823 (.A(net825),
    .X(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout824 (.A(net825),
    .X(net824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout825 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .X(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout826 (.A(net1042),
    .X(net826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout827 (.A(net828),
    .X(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout828 (.A(net268),
    .X(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout829 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .X(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout830 (.A(net832),
    .X(net830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout831 (.A(net832),
    .X(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout832 (.A(net1046),
    .X(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout833 (.A(net1044),
    .X(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout834 (.A(net977),
    .X(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout835 (.A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .X(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout836 (.A(net986),
    .X(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout837 (.A(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .X(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout838 (.A(\u_usb_cdc.u_sie.phy_state_q[9] ),
    .X(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout839 (.A(\u_usb_cdc.u_sie.phy_state_q[9] ),
    .X(net839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout840 (.A(net841),
    .X(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout841 (.A(net1017),
    .X(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout842 (.A(net843),
    .X(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout843 (.A(net1026),
    .X(net843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout844 (.A(net921),
    .X(net844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout845 (.A(net846),
    .X(net845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout846 (.A(net1035),
    .X(net846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout847 (.A(net848),
    .X(net847),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout848 (.A(net1047),
    .X(net848),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout849 (.A(net969),
    .X(net849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout850 (.A(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .X(net850),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout851 (.A(net513),
    .X(net851),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(usb_dn_rx_i),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(usb_dp_rx_i),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(usb_dn_en_o),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(usb_dn_tx_o),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(usb_dp_en_o),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(usb_dp_tx_o),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(usb_dp_up_o),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_usb_cdc_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net32));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_0_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_1_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk_regs (.A(clknet_3_2__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk_regs (.A(clknet_3_3__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk_regs (.A(clknet_3_7__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk_regs (.A(clknet_3_6__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_40_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_41_clk_regs (.A(clknet_3_5__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_42_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_43_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_44_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_45_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_46_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_47_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_47_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_48_clk_regs (.A(clknet_3_4__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_49_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_50_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_51_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_52_clk_regs (.A(clknet_3_1__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_53_clk_regs (.A(clknet_3_0__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload0 (.A(clknet_3_0__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_3_7__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload2 (.VDD(VPWR),
    .A(clknet_leaf_38_clk_regs),
    .VSS(VGND));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_21_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload4 (.VDD(VPWR),
    .A(clknet_leaf_34_clk_regs),
    .VSS(VGND));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_27_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_usb_cdc.rstn_sq[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_usb_cdc.clk_cnt_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold8 (.A(_1331_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0247_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_usb_cdc.u_sie.out_toggle_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0068_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0390_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0126_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_usb_cdc.clk_cnt_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0123_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0124_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0177_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0153_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0129_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0104_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0125_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0093_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0094_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0132_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0091_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_usb_cdc.u_sie.in_zlp_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0425_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0134_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0131_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0127_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0147_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0103_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0130_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0214_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0224_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0176_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0098_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_usb_cdc.u_sie.out_eop_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0360_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0149_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0179_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0120_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0182_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold74 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0128_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0095_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0106_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0150_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0202_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0210_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0232_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0096_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold90 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0151_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0135_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold94 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0154_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold96 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0152_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0050_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold100 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0200_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold103 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0208_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold105 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0230_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold107 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0138_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0231_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0117_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_usb_cdc.u_sie.delay_cnt_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0318_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold115 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0115_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0197_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0212_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold121 (.A(\u_usb_cdc.u_sie.in_zlp_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0426_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0237_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0100_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0238_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold129 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0191_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0052_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0209_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold134 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0122_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_usb_cdc.u_ctrl_endp.dev_state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold137 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0201_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0101_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold142 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0203_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_usb_cdc.u_sie.rx_data[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0401_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0204_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold148 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[67] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0092_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0121_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0118_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0148_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0175_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0119_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold164 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[66] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0233_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0362_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold168 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold171 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0207_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0167_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0116_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0097_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0181_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0223_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0236_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_usb_cdc.u_sie.rx_data[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0405_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0211_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_usb_cdc.u_sie.rx_data[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0403_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold191 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0213_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_usb_cdc.u_sie.rx_data[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0406_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0105_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0136_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0137_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold201 (.A(net24),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0248_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold203 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[38] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0205_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0102_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold207 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0099_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold209 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0133_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold212 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0173_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold214 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0199_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold216 (.A(net21),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0245_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold218 (.A(\u_usb_cdc.u_sie.addr_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold219 (.A(_1006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0072_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold221 (.A(net26),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0250_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_usb_cdc.u_sie.rx_data[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0404_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold225 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0180_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold227 (.A(\u_usb_cdc.u_sie.rx_data[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0408_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold229 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0196_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold231 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0387_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold233 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0225_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0178_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold237 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0195_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0376_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_usb_cdc.u_sie.rx_data[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold242 (.A(_1814_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold243 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0172_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold245 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0169_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold247 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0193_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0414_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold251 (.A(net25),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0249_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold253 (.A(net20),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0244_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold255 (.A(\u_usb_cdc.sie_out_data[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0054_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0073_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold258 (.A(\u_usb_cdc.u_sie.phy_state_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold260 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold261 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold262 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_err_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0944_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0058_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0418_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold267 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0365_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold269 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0361_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold271 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold273 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold274 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0215_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold276 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0383_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold278 (.A(\u_usb_cdc.u_sie.in_byte_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0321_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold280 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0228_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold282 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0185_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_usb_cdc.u_sie.in_byte_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0319_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0364_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold288 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0186_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold290 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold291 (.A(_1191_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0190_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold293 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0372_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0366_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold297 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0380_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold299 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold300 (.A(_1224_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0216_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold302 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0189_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold304 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[51] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold305 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0374_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold307 (.A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0422_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold309 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold310 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold311 (.A(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0316_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold313 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0415_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold315 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold316 (.A(_1187_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0188_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold318 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0370_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold320 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0166_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold322 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold323 (.A(_1751_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0371_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0037_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold327 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0198_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold329 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0229_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold331 (.A(\u_usb_cdc.u_sie.u_phy_rx.se0_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0421_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold333 (.A(\u_usb_cdc.u_sie.in_byte_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0320_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold335 (.A(\u_usb_cdc.u_sie.in_toggle_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0998_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0071_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold338 (.A(\u_usb_cdc.u_sie.addr_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0311_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold340 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0413_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold342 (.A(\u_usb_cdc.u_sie.addr_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0308_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold344 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0375_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold346 (.A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0423_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold348 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0379_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_usb_cdc.u_sie.u_phy_rx.state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0919_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0033_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold353 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold354 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold355 (.A(_1177_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0183_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold357 (.A(\u_usb_cdc.u_sie.in_byte_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0322_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold359 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0220_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold361 (.A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0424_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold363 (.A(\u_usb_cdc.u_sie.in_toggle_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0069_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold365 (.A(\u_usb_cdc.u_sie.addr_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold366 (.A(\u_usb_cdc.u_sie.addr_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0312_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold368 (.A(\u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold370 (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold371 (.A(_1471_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0314_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold373 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0217_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold375 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold376 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0165_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold378 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0363_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold380 (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold381 (.A(_1800_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0389_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold383 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0221_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold385 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0277_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold387 (.A(\u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold388 (.A(_1479_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0317_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold390 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0086_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold392 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0281_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold394 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0381_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold396 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold397 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold398 (.A(_1179_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0184_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold400 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0087_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold402 (.A(net22),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold403 (.A(_1313_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0246_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold405 (.A(\u_usb_cdc.u_sie.addr_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold406 (.A(\u_usb_cdc.u_sie.addr_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold407 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_valid_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0045_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold409 (.A(\u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold410 (.A(_1811_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0398_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold412 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0088_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold414 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0378_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold417 (.A(_1882_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold418 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0083_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold420 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0144_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold422 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0392_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold424 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold426 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0141_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold428 (.A(\u_usb_cdc.u_ctrl_endp.state_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0015_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold430 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0280_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold432 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0143_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold434 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0146_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold436 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold437 (.A(_0145_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0060_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0420_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold440 (.A(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold442 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold443 (.A(\u_usb_cdc.u_sie.out_toggle_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0067_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold445 (.A(\u_usb_cdc.u_sie.data_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0055_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold447 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0085_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold449 (.A(\u_usb_cdc.u_ctrl_endp.class_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0286_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold451 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold452 (.A(_1876_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold453 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0367_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold455 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold456 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold457 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold458 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0945_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold461 (.A(\u_usb_cdc.u_sie.phy_state_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold463 (.A(\u_usb_cdc.u_sie.rx_data[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold464 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0139_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold466 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0114_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold468 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0108_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold470 (.A(\u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold472 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0107_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold474 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0140_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold476 (.A(\u_usb_cdc.u_sie.data_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold477 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0112_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold479 (.A(\u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0001_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold481 (.A(\u_usb_cdc.u_sie.phy_state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold483 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0089_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold485 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0110_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold487 (.A(\u_usb_cdc.u_sie.crc16_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0323_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold489 (.A(\u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold490 (.A(_1812_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0399_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold492 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0111_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold494 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0109_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold496 (.A(\u_usb_cdc.u_sie.crc16_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0336_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0062_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold500 (.A(\u_usb_cdc.out_valid_o [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold502 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0265_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold504 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0074_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold506 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0084_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold508 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold509 (.A(_1907_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold510 (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold511 (.A(_1809_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold512 (.A(_0396_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold513 (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold514 (.A(_1810_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold515 (.A(_0397_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold516 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold517 (.A(\u_usb_cdc.u_sie.data_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0866_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold519 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0301_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold521 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0294_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold523 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold524 (.A(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold525 (.A(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0920_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold527 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0113_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold529 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0893_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold532 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0164_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold534 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold535 (.A(\u_usb_cdc.u_sie.crc16_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold536 (.A(_0333_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold537 (.A(\u_usb_cdc.u_sie.in_toggle_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0993_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold539 (.A(_0070_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold540 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold541 (.A(_0155_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold542 (.A(\u_usb_cdc.addr[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold543 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0156_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold545 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0290_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold547 (.A(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0003_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold549 (.A(\u_usb_cdc.addr[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold550 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold552 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold553 (.A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold554 (.A(_2029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold555 (.A(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold557 (.A(\u_usb_cdc.u_sie.rx_err ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0393_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold559 (.A(\u_usb_cdc.addr[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold560 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold561 (.A(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold562 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold563 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold564 (.A(_0157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold565 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold566 (.A(net31),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold567 (.A(_1820_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold568 (.A(_0409_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_usb_cdc.u_sie.crc16_q[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0332_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold571 (.A(\u_usb_cdc.u_sie.crc16_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold572 (.A(_0330_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold573 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold574 (.A(_0240_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold575 (.A(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold576 (.A(_0002_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold577 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold578 (.A(\u_usb_cdc.addr[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold579 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0291_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold581 (.A(\u_usb_cdc.addr[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold582 (.A(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold583 (.A(\u_usb_cdc.u_sie.crc16_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold584 (.A(_0334_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold585 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold586 (.A(\u_usb_cdc.addr[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold587 (.A(\u_usb_cdc.u_sie.crc16_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0329_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold589 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0293_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold591 (.A(\u_usb_cdc.u_sie.crc16_q[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold592 (.A(\u_usb_cdc.u_sie.pid_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold593 (.A(_0355_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold594 (.A(\u_usb_cdc.u_sie.crc16_q[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0335_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold596 (.A(\u_usb_cdc.u_sie.crc16_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold597 (.A(_0331_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold598 (.A(\u_usb_cdc.bus_reset ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold599 (.A(_1803_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0391_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold601 (.A(\u_usb_cdc.u_sie.crc16_q[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold602 (.A(\u_usb_cdc.u_sie.phy_state_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold603 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold604 (.A(\u_usb_cdc.addr[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold605 (.A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold606 (.A(_0928_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold607 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold608 (.A(_0289_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold609 (.A(\u_usb_cdc.u_sie.crc16_q[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold610 (.A(\u_usb_cdc.u_sie.u_phy_rx.state_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold611 (.A(_0035_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold612 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold613 (.A(\u_usb_cdc.u_sie.crc16_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold614 (.A(\u_usb_cdc.in_ready_o [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold615 (.A(\u_usb_cdc.u_sie.rx_valid ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold616 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold617 (.A(_0252_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold618 (.A(_0059_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0048_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold620 (.A(_0061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold621 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold622 (.A(_0253_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold623 (.A(\u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold624 (.A(_0004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold625 (.A(\u_usb_cdc.u_sie.pid_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold626 (.A(_0356_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold627 (.A(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0836_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold630 (.A(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold631 (.A(_0017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold632 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold633 (.A(_0254_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold634 (.A(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold635 (.A(_0285_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold636 (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold637 (.A(_0313_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold638 (.A(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold639 (.A(_0008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold640 (.A(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold642 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold643 (.A(_1740_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold644 (.A(_1741_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold645 (.A(_0368_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold646 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold647 (.A(_0258_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold648 (.A(\u_usb_cdc.u_sie.crc16_q[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold649 (.A(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold650 (.A(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold651 (.A(_0013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold652 (.A(\u_usb_cdc.endp[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold653 (.A(\u_usb_cdc.endp[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold654 (.A(\u_usb_cdc.u_sie.crc16_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold655 (.A(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold656 (.A(_0009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold657 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold658 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold659 (.A(_0159_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold660 (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold661 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold662 (.A(_0262_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold663 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold664 (.A(_0373_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold665 (.A(\u_usb_cdc.u_sie.data_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold666 (.A(net19),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold667 (.A(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold668 (.A(_0580_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold669 (.A(_0581_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold670 (.A(\u_usb_cdc.u_sie.data_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold671 (.A(_0051_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold672 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold673 (.A(\u_usb_cdc.u_sie.data_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold674 (.A(\u_usb_cdc.endp[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold675 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold676 (.A(\u_usb_cdc.endp[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold677 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold678 (.A(\u_usb_cdc.u_sie.data_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold679 (.A(\u_usb_cdc.u_sie.pid_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0357_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold681 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold682 (.A(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold683 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold684 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold685 (.A(_0251_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold686 (.A(\u_usb_cdc.u_sie.data_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold687 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold688 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold689 (.A(_0030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold690 (.A(_0060_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold691 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold692 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold693 (.A(\u_usb_cdc.sie_out_data[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold694 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold695 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold696 (.A(_1377_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold697 (.A(_0260_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold698 (.A(\u_usb_cdc.u_sie.phy_state_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold699 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold700 (.A(\u_usb_cdc.sie_out_data[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold701 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold702 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold703 (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold704 (.A(_0064_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold705 (.A(\u_usb_cdc.sie_out_data[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold706 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold707 (.A(\u_usb_cdc.u_sie.phy_state_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold708 (.A(_0875_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold709 (.A(\u_usb_cdc.u_sie.pid_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold710 (.A(_0358_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold711 (.A(\u_usb_cdc.ctrl_stall ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold712 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold713 (.A(_0257_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold714 (.A(\u_usb_cdc.sie_out_data[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold715 (.A(\u_usb_cdc.sie_in_req ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold716 (.A(\u_usb_cdc.u_sie.phy_state_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold717 (.A(_0879_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold718 (.A(\u_usb_cdc.sie_in_data_ack ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold719 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0056_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold721 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold722 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold723 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold724 (.A(\u_usb_cdc.sie_out_err ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold725 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold726 (.A(\u_usb_cdc.sie_out_data[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold727 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold728 (.A(\u_usb_cdc.u_sie.phy_state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold729 (.A(\u_usb_cdc.rstn ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold730 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold731 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold732 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold733 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold734 (.A(\u_usb_cdc.u_sie.pid_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold735 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1054));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net32;
 assign uio_oe[1] = net33;
 assign uio_oe[2] = net34;
 assign uio_oe[3] = net39;
 assign uio_oe[4] = net40;
 assign uio_oe[5] = net41;
 assign uio_oe[6] = net42;
 assign uio_oe[7] = net43;
 assign uio_out[0] = net35;
 assign uio_out[1] = net36;
 assign uio_out[2] = net37;
endmodule
