module heichips25_usb_cdc (clk,
    ena,
    rst_n,
    usb_dn_en_o,
    usb_dn_rx_i,
    usb_dn_tx_o,
    usb_dp_en_o,
    usb_dp_rx_i,
    usb_dp_tx_o,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 output usb_dn_en_o;
 input usb_dn_rx_i;
 output usb_dn_tx_o;
 output usb_dp_en_o;
 input usb_dp_rx_i;
 output usb_dp_tx_o;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire clknet_leaf_0_clk;
 wire \u_usb_cdc.addr[0] ;
 wire \u_usb_cdc.addr[1] ;
 wire \u_usb_cdc.addr[2] ;
 wire \u_usb_cdc.addr[3] ;
 wire \u_usb_cdc.addr[4] ;
 wire \u_usb_cdc.addr[5] ;
 wire \u_usb_cdc.addr[6] ;
 wire \u_usb_cdc.bus_reset ;
 wire \u_usb_cdc.clk_cnt_q[0] ;
 wire \u_usb_cdc.clk_cnt_q[1] ;
 wire \u_usb_cdc.clk_gate_q ;
 wire \u_usb_cdc.configured_o ;
 wire \u_usb_cdc.ctrl_stall ;
 wire \u_usb_cdc.dp_pu_o ;
 wire \u_usb_cdc.endp[0] ;
 wire \u_usb_cdc.endp[1] ;
 wire \u_usb_cdc.endp[2] ;
 wire \u_usb_cdc.endp[3] ;
 wire \u_usb_cdc.rstn ;
 wire \u_usb_cdc.rstn_sq[1] ;
 wire \u_usb_cdc.sie_in_data_ack ;
 wire \u_usb_cdc.sie_in_req ;
 wire \u_usb_cdc.sie_out_data[0] ;
 wire \u_usb_cdc.sie_out_data[1] ;
 wire \u_usb_cdc.sie_out_data[2] ;
 wire \u_usb_cdc.sie_out_data[3] ;
 wire \u_usb_cdc.sie_out_data[4] ;
 wire \u_usb_cdc.sie_out_data[5] ;
 wire \u_usb_cdc.sie_out_data[6] ;
 wire \u_usb_cdc.sie_out_data[7] ;
 wire \u_usb_cdc.sie_out_err ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[63] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[71] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[11] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[14] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[18] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[23] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[26] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[28] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[29] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[31] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[35] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[38] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[51] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[54] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[59] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[62] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[64] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[65] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[66] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[67] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[68] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[69] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[6] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[70] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[71] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ;
 wire \u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[0] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[1] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[2] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[3] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[4] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[5] ;
 wire \u_usb_cdc.u_ctrl_endp.addr_dd[6] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.class_q ;
 wire \u_usb_cdc.u_ctrl_endp.dev_state_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ;
 wire \u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.endp_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.in_dir_q ;
 wire \u_usb_cdc.u_ctrl_endp.in_endp_q ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[4] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.max_length_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.rec_q[0] ;
 wire \u_usb_cdc.u_ctrl_endp.rec_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[10] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[11] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[4] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[7] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[8] ;
 wire \u_usb_cdc.u_ctrl_endp.req_q[9] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[1] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[2] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[3] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[5] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[6] ;
 wire \u_usb_cdc.u_ctrl_endp.state_q[7] ;
 wire \u_usb_cdc.u_sie.addr_q[0] ;
 wire \u_usb_cdc.u_sie.addr_q[1] ;
 wire \u_usb_cdc.u_sie.addr_q[2] ;
 wire \u_usb_cdc.u_sie.addr_q[3] ;
 wire \u_usb_cdc.u_sie.addr_q[4] ;
 wire \u_usb_cdc.u_sie.addr_q[5] ;
 wire \u_usb_cdc.u_sie.addr_q[6] ;
 wire \u_usb_cdc.u_sie.crc16_q[0] ;
 wire \u_usb_cdc.u_sie.crc16_q[10] ;
 wire \u_usb_cdc.u_sie.crc16_q[11] ;
 wire \u_usb_cdc.u_sie.crc16_q[12] ;
 wire \u_usb_cdc.u_sie.crc16_q[13] ;
 wire \u_usb_cdc.u_sie.crc16_q[14] ;
 wire \u_usb_cdc.u_sie.crc16_q[15] ;
 wire \u_usb_cdc.u_sie.crc16_q[1] ;
 wire \u_usb_cdc.u_sie.crc16_q[2] ;
 wire \u_usb_cdc.u_sie.crc16_q[3] ;
 wire \u_usb_cdc.u_sie.crc16_q[4] ;
 wire \u_usb_cdc.u_sie.crc16_q[5] ;
 wire \u_usb_cdc.u_sie.crc16_q[6] ;
 wire \u_usb_cdc.u_sie.crc16_q[7] ;
 wire \u_usb_cdc.u_sie.crc16_q[8] ;
 wire \u_usb_cdc.u_sie.crc16_q[9] ;
 wire \u_usb_cdc.u_sie.data_q[0] ;
 wire \u_usb_cdc.u_sie.data_q[1] ;
 wire \u_usb_cdc.u_sie.data_q[2] ;
 wire \u_usb_cdc.u_sie.data_q[3] ;
 wire \u_usb_cdc.u_sie.data_q[4] ;
 wire \u_usb_cdc.u_sie.data_q[5] ;
 wire \u_usb_cdc.u_sie.data_q[6] ;
 wire \u_usb_cdc.u_sie.data_q[7] ;
 wire \u_usb_cdc.u_sie.delay_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.delay_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.delay_cnt_q[2] ;
 wire \u_usb_cdc.u_sie.in_byte_q[0] ;
 wire \u_usb_cdc.u_sie.in_byte_q[1] ;
 wire \u_usb_cdc.u_sie.in_byte_q[2] ;
 wire \u_usb_cdc.u_sie.in_byte_q[3] ;
 wire \u_usb_cdc.u_sie.in_toggle_q[0] ;
 wire \u_usb_cdc.u_sie.in_toggle_q[1] ;
 wire \u_usb_cdc.u_sie.in_toggle_q[2] ;
 wire \u_usb_cdc.u_sie.in_zlp_q[0] ;
 wire \u_usb_cdc.u_sie.in_zlp_q[1] ;
 wire \u_usb_cdc.u_sie.out_eop_q ;
 wire \u_usb_cdc.u_sie.out_toggle_q[0] ;
 wire \u_usb_cdc.u_sie.out_toggle_q[1] ;
 wire \u_usb_cdc.u_sie.phy_state_q[10] ;
 wire \u_usb_cdc.u_sie.phy_state_q[11] ;
 wire \u_usb_cdc.u_sie.phy_state_q[1] ;
 wire \u_usb_cdc.u_sie.phy_state_q[2] ;
 wire \u_usb_cdc.u_sie.phy_state_q[3] ;
 wire \u_usb_cdc.u_sie.phy_state_q[4] ;
 wire \u_usb_cdc.u_sie.phy_state_q[5] ;
 wire \u_usb_cdc.u_sie.phy_state_q[6] ;
 wire \u_usb_cdc.u_sie.phy_state_q[7] ;
 wire \u_usb_cdc.u_sie.phy_state_q[8] ;
 wire \u_usb_cdc.u_sie.phy_state_q[9] ;
 wire \u_usb_cdc.u_sie.pid_q[0] ;
 wire \u_usb_cdc.u_sie.pid_q[1] ;
 wire \u_usb_cdc.u_sie.pid_q[2] ;
 wire \u_usb_cdc.u_sie.pid_q[3] ;
 wire \u_usb_cdc.u_sie.rx_data[0] ;
 wire \u_usb_cdc.u_sie.rx_data[1] ;
 wire \u_usb_cdc.u_sie.rx_data[2] ;
 wire \u_usb_cdc.u_sie.rx_data[3] ;
 wire \u_usb_cdc.u_sie.rx_data[4] ;
 wire \u_usb_cdc.u_sie.rx_data[5] ;
 wire \u_usb_cdc.u_sie.rx_data[6] ;
 wire \u_usb_cdc.u_sie.rx_data[7] ;
 wire \u_usb_cdc.u_sie.rx_err ;
 wire \u_usb_cdc.u_sie.rx_valid ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_en_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_eop_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_err_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.rx_valid_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.se0_q ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[5] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.state_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.state_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.state_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[3] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[4] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[5] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.data_q[6] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ;
 wire \u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net42;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net41;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire [0:0] \u_usb_cdc.bulk_out_nak ;
 wire [0:0] \u_usb_cdc.in_ready_o ;
 wire [0:0] \u_usb_cdc.out_valid_o ;

 sg13g2_inv_1 _2014_ (.Y(_1893_),
    .A(net308));
 sg13g2_inv_4 _2015_ (.A(net761),
    .Y(_1894_));
 sg13g2_inv_4 _2016_ (.A(net757),
    .Y(_1895_));
 sg13g2_inv_1 _2017_ (.Y(_1896_),
    .A(net755));
 sg13g2_inv_1 _2018_ (.Y(_1897_),
    .A(net756));
 sg13g2_inv_8 _2019_ (.Y(_1898_),
    .A(net753));
 sg13g2_inv_4 _2020_ (.A(net754),
    .Y(_1899_));
 sg13g2_inv_4 _2021_ (.A(net751),
    .Y(_1900_));
 sg13g2_inv_8 _2022_ (.Y(_1901_),
    .A(net752));
 sg13g2_inv_1 _2023_ (.Y(_1902_),
    .A(net745));
 sg13g2_inv_1 _2024_ (.Y(_1903_),
    .A(net833));
 sg13g2_inv_4 _2025_ (.A(net747),
    .Y(_1904_));
 sg13g2_inv_1 _2026_ (.Y(_1905_),
    .A(net884));
 sg13g2_inv_2 _2027_ (.Y(_1906_),
    .A(net767));
 sg13g2_inv_1 _2028_ (.Y(_1907_),
    .A(net958));
 sg13g2_inv_1 _2029_ (.Y(_1908_),
    .A(net964));
 sg13g2_inv_1 _2030_ (.Y(_1909_),
    .A(net1034));
 sg13g2_inv_2 _2031_ (.Y(_1910_),
    .A(net835));
 sg13g2_inv_1 _2032_ (.Y(_1911_),
    .A(net829));
 sg13g2_inv_2 _2033_ (.Y(_1912_),
    .A(net803));
 sg13g2_inv_4 _2034_ (.A(net989),
    .Y(_1913_));
 sg13g2_inv_2 _2035_ (.Y(_1914_),
    .A(net788));
 sg13g2_inv_4 _2036_ (.A(net786),
    .Y(_1915_));
 sg13g2_inv_1 _2037_ (.Y(_1916_),
    .A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ));
 sg13g2_inv_2 _2038_ (.Y(_1917_),
    .A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ));
 sg13g2_inv_1 _2039_ (.Y(_1918_),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[2] ));
 sg13g2_inv_1 _2040_ (.Y(_1919_),
    .A(net866));
 sg13g2_inv_1 _2041_ (.Y(_1920_),
    .A(net1003));
 sg13g2_inv_1 _2042_ (.Y(_1921_),
    .A(net460));
 sg13g2_inv_1 _2043_ (.Y(_1922_),
    .A(\u_usb_cdc.u_sie.pid_q[0] ));
 sg13g2_inv_1 _2044_ (.Y(_1923_),
    .A(\u_usb_cdc.u_sie.pid_q[1] ));
 sg13g2_inv_2 _2045_ (.Y(_1924_),
    .A(\u_usb_cdc.u_sie.pid_q[2] ));
 sg13g2_inv_2 _2046_ (.Y(_1925_),
    .A(\u_usb_cdc.u_sie.pid_q[3] ));
 sg13g2_inv_2 _2047_ (.Y(_1926_),
    .A(net920));
 sg13g2_inv_2 _2048_ (.Y(_1927_),
    .A(net910));
 sg13g2_inv_1 _2049_ (.Y(_1928_),
    .A(\u_usb_cdc.u_ctrl_endp.in_dir_q ));
 sg13g2_inv_1 _2050_ (.Y(_1929_),
    .A(net741));
 sg13g2_inv_1 _2051_ (.Y(_1930_),
    .A(net868));
 sg13g2_inv_1 _2052_ (.Y(_1931_),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[6] ));
 sg13g2_inv_2 _2053_ (.Y(_1932_),
    .A(net842));
 sg13g2_inv_1 _2054_ (.Y(_1933_),
    .A(net949));
 sg13g2_inv_2 _2055_ (.Y(_1934_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ));
 sg13g2_inv_4 _2056_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .Y(_1935_));
 sg13g2_inv_1 _2057_ (.Y(_1936_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ));
 sg13g2_inv_2 _2058_ (.Y(_1937_),
    .A(net935));
 sg13g2_inv_1 _2059_ (.Y(_1938_),
    .A(net915));
 sg13g2_inv_1 _2060_ (.Y(_1939_),
    .A(\u_usb_cdc.u_sie.crc16_q[14] ));
 sg13g2_inv_1 _2061_ (.Y(_1940_),
    .A(\u_usb_cdc.u_sie.crc16_q[13] ));
 sg13g2_inv_1 _2062_ (.Y(_1941_),
    .A(\u_usb_cdc.u_sie.crc16_q[12] ));
 sg13g2_inv_1 _2063_ (.Y(_1942_),
    .A(\u_usb_cdc.u_sie.crc16_q[11] ));
 sg13g2_inv_1 _2064_ (.Y(_1943_),
    .A(net444));
 sg13g2_inv_1 _2065_ (.Y(_1944_),
    .A(net540));
 sg13g2_inv_1 _2066_ (.Y(_1945_),
    .A(net881));
 sg13g2_inv_2 _2067_ (.Y(_1946_),
    .A(net409));
 sg13g2_inv_1 _2068_ (.Y(_1947_),
    .A(net918));
 sg13g2_inv_2 _2069_ (.Y(_1948_),
    .A(net372));
 sg13g2_inv_1 _2070_ (.Y(_1949_),
    .A(net502));
 sg13g2_inv_2 _2071_ (.Y(_1950_),
    .A(net306));
 sg13g2_inv_2 _2072_ (.Y(_1951_),
    .A(net285));
 sg13g2_inv_2 _2073_ (.Y(_1952_),
    .A(net882));
 sg13g2_inv_2 _2074_ (.Y(_1953_),
    .A(net349));
 sg13g2_inv_1 _2075_ (.Y(_1954_),
    .A(\u_usb_cdc.addr[0] ));
 sg13g2_inv_1 _2076_ (.Y(_1955_),
    .A(net479));
 sg13g2_inv_1 _2077_ (.Y(_1956_),
    .A(net186));
 sg13g2_inv_1 _2078_ (.Y(_1957_),
    .A(net525));
 sg13g2_inv_1 _2079_ (.Y(_1958_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ));
 sg13g2_inv_1 _2080_ (.Y(_1959_),
    .A(net189));
 sg13g2_inv_1 _2081_ (.Y(_1960_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ));
 sg13g2_inv_1 _2082_ (.Y(_1961_),
    .A(net987));
 sg13g2_inv_1 _2083_ (.Y(_1962_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ));
 sg13g2_inv_2 _2084_ (.Y(_1963_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ));
 sg13g2_inv_2 _2085_ (.Y(_1964_),
    .A(net1069));
 sg13g2_inv_2 _2086_ (.Y(_1965_),
    .A(net826));
 sg13g2_inv_1 _2087_ (.Y(_0039_),
    .A(net48));
 sg13g2_inv_2 _2088_ (.Y(_1966_),
    .A(net310));
 sg13g2_inv_1 _2089_ (.Y(_1967_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ));
 sg13g2_inv_1 _2090_ (.Y(_1968_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ));
 sg13g2_inv_1 _2091_ (.Y(_1969_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ));
 sg13g2_inv_1 _2092_ (.Y(_1970_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ));
 sg13g2_inv_1 _2093_ (.Y(_1971_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ));
 sg13g2_inv_1 _2094_ (.Y(_1972_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ));
 sg13g2_inv_1 _2095_ (.Y(_1973_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ));
 sg13g2_inv_1 _2096_ (.Y(_1974_),
    .A(net337));
 sg13g2_inv_2 _2097_ (.Y(_1975_),
    .A(net979));
 sg13g2_inv_1 _2098_ (.Y(_1976_),
    .A(net265));
 sg13g2_inv_1 _2099_ (.Y(_1977_),
    .A(net466));
 sg13g2_inv_1 _2100_ (.Y(_1978_),
    .A(net102));
 sg13g2_inv_1 _2101_ (.Y(_1979_),
    .A(net180));
 sg13g2_inv_1 _2102_ (.Y(_1980_),
    .A(net244));
 sg13g2_inv_1 _2103_ (.Y(_1981_),
    .A(net287));
 sg13g2_inv_1 _2104_ (.Y(_1982_),
    .A(net860));
 sg13g2_inv_1 _2105_ (.Y(_1983_),
    .A(net136));
 sg13g2_inv_1 _2106_ (.Y(_1984_),
    .A(net382));
 sg13g2_or2_1 _2107_ (.X(_1985_),
    .B(\u_usb_cdc.endp[2] ),
    .A(\u_usb_cdc.endp[1] ));
 sg13g2_nor3_2 _2108_ (.A(\u_usb_cdc.endp[1] ),
    .B(\u_usb_cdc.endp[3] ),
    .C(\u_usb_cdc.endp[2] ),
    .Y(_1986_));
 sg13g2_nor2_1 _2109_ (.A(net767),
    .B(\u_usb_cdc.endp[2] ),
    .Y(_1987_));
 sg13g2_nor3_1 _2110_ (.A(net767),
    .B(\u_usb_cdc.endp[3] ),
    .C(\u_usb_cdc.endp[2] ),
    .Y(_1988_));
 sg13g2_nor2_2 _2111_ (.A(net706),
    .B(_1988_),
    .Y(_1989_));
 sg13g2_nor2b_1 _2112_ (.A(_1989_),
    .B_N(net839),
    .Y(_1990_));
 sg13g2_o21ai_1 _2113_ (.B1(net839),
    .Y(_1991_),
    .A1(net706),
    .A2(_1988_));
 sg13g2_nor4_1 _2114_ (.A(net838),
    .B(net834),
    .C(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .D(net831),
    .Y(_1992_));
 sg13g2_a21oi_2 _2115_ (.B1(net747),
    .Y(_1993_),
    .A2(_1992_),
    .A1(_1991_));
 sg13g2_a21o_2 _2116_ (.A2(_1992_),
    .A1(_1991_),
    .B1(net748),
    .X(_1994_));
 sg13g2_nand2_1 _2117_ (.Y(_1995_),
    .A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .B(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ));
 sg13g2_nor2_1 _2118_ (.A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_or2_1 _2119_ (.X(_1997_),
    .B(_1995_),
    .A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ));
 sg13g2_nor2_1 _2120_ (.A(net713),
    .B(_1996_),
    .Y(_1998_));
 sg13g2_nand2_2 _2121_ (.Y(_1999_),
    .A(net743),
    .B(_1997_));
 sg13g2_nand2_1 _2122_ (.Y(_2000_),
    .A(_1993_),
    .B(net623));
 sg13g2_nand2_1 _2123_ (.Y(_2001_),
    .A(net312),
    .B(net210));
 sg13g2_and3_2 _2124_ (.X(_2002_),
    .A(_0060_),
    .B(net312),
    .C(_0058_));
 sg13g2_nand3_1 _2125_ (.B(net312),
    .C(net210),
    .A(_0060_),
    .Y(_2003_));
 sg13g2_nor2_1 _2126_ (.A(_1993_),
    .B(_2003_),
    .Y(_2004_));
 sg13g2_nand2_1 _2127_ (.Y(_2005_),
    .A(_1994_),
    .B(net705));
 sg13g2_nand2_1 _2128_ (.Y(_2006_),
    .A(net931),
    .B(_2004_));
 sg13g2_o21ai_1 _2129_ (.B1(_2006_),
    .Y(_2007_),
    .A1(_1911_),
    .A2(_2003_));
 sg13g2_a22oi_1 _2130_ (.Y(_0066_),
    .B1(_2007_),
    .B2(net623),
    .A2(_2000_),
    .A1(_1984_));
 sg13g2_nand2_1 _2131_ (.Y(_0065_),
    .A(net712),
    .B(_1983_));
 sg13g2_nor2b_2 _2132_ (.A(net988),
    .B_N(net973),
    .Y(_2008_));
 sg13g2_nor2b_1 _2133_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .B_N(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .Y(_2009_));
 sg13g2_nor2_1 _2134_ (.A(_1934_),
    .B(net973),
    .Y(_2010_));
 sg13g2_nor2_1 _2135_ (.A(_1935_),
    .B(net913),
    .Y(_2011_));
 sg13g2_nor4_2 _2136_ (.A(_2008_),
    .B(_2009_),
    .C(_2010_),
    .Y(_2012_),
    .D(_2011_));
 sg13g2_nor2_2 _2137_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .Y(_0440_));
 sg13g2_nand2_2 _2138_ (.Y(_0441_),
    .A(_1934_),
    .B(_1935_));
 sg13g2_nor2_1 _2139_ (.A(_1934_),
    .B(_1935_),
    .Y(_0442_));
 sg13g2_nor3_2 _2140_ (.A(_2012_),
    .B(_0440_),
    .C(_0442_),
    .Y(_0443_));
 sg13g2_inv_1 _2141_ (.Y(_0444_),
    .A(_0443_));
 sg13g2_nor4_1 _2142_ (.A(_1935_),
    .B(net899),
    .C(net862),
    .D(net908),
    .Y(_0445_));
 sg13g2_nor2_1 _2143_ (.A(net428),
    .B(net527),
    .Y(_0446_));
 sg13g2_and4_1 _2144_ (.A(net360),
    .B(_1934_),
    .C(_0445_),
    .D(_0446_),
    .X(_0447_));
 sg13g2_nor2b_2 _2145_ (.A(net521),
    .B_N(net49),
    .Y(_0448_));
 sg13g2_nand2b_1 _2146_ (.Y(_0449_),
    .B(net49),
    .A_N(net521));
 sg13g2_nor2_2 _2147_ (.A(_1937_),
    .B(net703),
    .Y(_0450_));
 sg13g2_nand2_1 _2148_ (.Y(_0451_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .B(_0450_));
 sg13g2_nor3_1 _2149_ (.A(_0443_),
    .B(_0447_),
    .C(_0451_),
    .Y(_0452_));
 sg13g2_nand2_1 _2150_ (.Y(_0453_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(_1935_));
 sg13g2_and4_1 _2151_ (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .B(_1935_),
    .C(net257),
    .D(net635),
    .X(_0454_));
 sg13g2_nand2_1 _2152_ (.Y(_0455_),
    .A(_2008_),
    .B(_2011_));
 sg13g2_a21oi_1 _2153_ (.A1(_2008_),
    .A2(_2011_),
    .Y(_0456_),
    .B1(net351));
 sg13g2_a22oi_1 _2154_ (.Y(_0457_),
    .B1(net635),
    .B2(_1958_),
    .A2(net703),
    .A1(net351));
 sg13g2_nor4_1 _2155_ (.A(_0452_),
    .B(_0454_),
    .C(net352),
    .D(_0457_),
    .Y(_0064_));
 sg13g2_xnor2_1 _2156_ (.Y(_0458_),
    .A(net753),
    .B(\u_usb_cdc.addr[5] ));
 sg13g2_xnor2_1 _2157_ (.Y(_0459_),
    .A(net752),
    .B(\u_usb_cdc.addr[6] ));
 sg13g2_xor2_1 _2158_ (.B(\u_usb_cdc.addr[1] ),
    .A(net758),
    .X(_0460_));
 sg13g2_xor2_1 _2159_ (.B(\u_usb_cdc.addr[4] ),
    .A(net754),
    .X(_0461_));
 sg13g2_xor2_1 _2160_ (.B(\u_usb_cdc.addr[0] ),
    .A(net760),
    .X(_0462_));
 sg13g2_xnor2_1 _2161_ (.Y(_0463_),
    .A(net755),
    .B(\u_usb_cdc.addr[3] ));
 sg13g2_xor2_1 _2162_ (.B(\u_usb_cdc.addr[2] ),
    .A(net756),
    .X(_0464_));
 sg13g2_nor4_1 _2163_ (.A(_0460_),
    .B(_0461_),
    .C(_0462_),
    .D(_0464_),
    .Y(_0465_));
 sg13g2_nand4_1 _2164_ (.B(_0459_),
    .C(_0463_),
    .A(_0458_),
    .Y(_0466_),
    .D(_0465_));
 sg13g2_nor2_1 _2165_ (.A(_1922_),
    .B(\u_usb_cdc.u_sie.pid_q[1] ),
    .Y(_0467_));
 sg13g2_nand2_1 _2166_ (.Y(_0468_),
    .A(net1018),
    .B(_0467_));
 sg13g2_or3_1 _2167_ (.A(net1009),
    .B(_0466_),
    .C(_0468_),
    .X(_0469_));
 sg13g2_xor2_1 _2168_ (.B(net754),
    .A(net758),
    .X(_0470_));
 sg13g2_xnor2_1 _2169_ (.Y(_0471_),
    .A(net756),
    .B(net751));
 sg13g2_xnor2_1 _2170_ (.Y(_0472_),
    .A(_0470_),
    .B(_0471_));
 sg13g2_xnor2_1 _2171_ (.Y(_0473_),
    .A(\u_usb_cdc.sie_out_data[2] ),
    .B(net753));
 sg13g2_xnor2_1 _2172_ (.Y(_0474_),
    .A(\u_usb_cdc.sie_out_data[0] ),
    .B(net762));
 sg13g2_xnor2_1 _2173_ (.Y(_0475_),
    .A(_0473_),
    .B(_0474_));
 sg13g2_xnor2_1 _2174_ (.Y(_0476_),
    .A(_0472_),
    .B(_0475_));
 sg13g2_xnor2_1 _2175_ (.Y(_0477_),
    .A(\u_usb_cdc.u_sie.data_q[7] ),
    .B(_0476_));
 sg13g2_nand2_1 _2176_ (.Y(_0478_),
    .A(net760),
    .B(net757));
 sg13g2_nor2_1 _2177_ (.A(net760),
    .B(net757),
    .Y(_0479_));
 sg13g2_nand2_2 _2178_ (.Y(_0480_),
    .A(net721),
    .B(net757));
 sg13g2_xor2_1 _2179_ (.B(net758),
    .A(net761),
    .X(_0481_));
 sg13g2_xnor2_1 _2180_ (.Y(_0482_),
    .A(\u_usb_cdc.sie_out_data[3] ),
    .B(net752));
 sg13g2_xnor2_1 _2181_ (.Y(_0483_),
    .A(_0481_),
    .B(_0482_));
 sg13g2_xnor2_1 _2182_ (.Y(_0484_),
    .A(net764),
    .B(_0470_));
 sg13g2_xnor2_1 _2183_ (.Y(_0485_),
    .A(_0483_),
    .B(_0484_));
 sg13g2_xor2_1 _2184_ (.B(_0472_),
    .A(\u_usb_cdc.u_sie.data_q[4] ),
    .X(_0486_));
 sg13g2_mux2_1 _2185_ (.A0(_0486_),
    .A1(_0485_),
    .S(\u_usb_cdc.u_sie.data_q[6] ),
    .X(_0487_));
 sg13g2_xnor2_1 _2186_ (.Y(_0488_),
    .A(\u_usb_cdc.sie_out_data[3] ),
    .B(net766));
 sg13g2_xnor2_1 _2187_ (.Y(_0489_),
    .A(_0473_),
    .B(_0488_));
 sg13g2_xor2_1 _2188_ (.B(_0483_),
    .A(\u_usb_cdc.u_sie.data_q[3] ),
    .X(_0490_));
 sg13g2_a22oi_1 _2189_ (.Y(_0491_),
    .B1(_0489_),
    .B2(_0490_),
    .A2(_0486_),
    .A1(_0485_));
 sg13g2_xor2_1 _2190_ (.B(_0476_),
    .A(\u_usb_cdc.u_sie.data_q[5] ),
    .X(_0492_));
 sg13g2_mux2_1 _2191_ (.A0(_0489_),
    .A1(_0490_),
    .S(_0492_),
    .X(_0493_));
 sg13g2_and4_1 _2192_ (.A(_0477_),
    .B(_0487_),
    .C(_0491_),
    .D(_0493_),
    .X(_0494_));
 sg13g2_nand2_1 _2193_ (.Y(_0495_),
    .A(\u_usb_cdc.u_sie.pid_q[2] ),
    .B(_1925_));
 sg13g2_nand3_1 _2194_ (.B(_1925_),
    .C(_0467_),
    .A(\u_usb_cdc.u_sie.pid_q[2] ),
    .Y(_0496_));
 sg13g2_inv_1 _2195_ (.Y(_0497_),
    .A(_0496_));
 sg13g2_nand2_1 _2196_ (.Y(_0498_),
    .A(_0494_),
    .B(_0496_));
 sg13g2_o21ai_1 _2197_ (.B1(net832),
    .Y(_0499_),
    .A1(_0469_),
    .A2(_0498_));
 sg13g2_xor2_1 _2198_ (.B(\u_usb_cdc.u_sie.data_q[7] ),
    .A(net881),
    .X(_0500_));
 sg13g2_xor2_1 _2199_ (.B(\u_usb_cdc.u_sie.data_q[6] ),
    .A(net540),
    .X(_0501_));
 sg13g2_xor2_1 _2200_ (.B(\u_usb_cdc.u_sie.data_q[5] ),
    .A(net444),
    .X(_0502_));
 sg13g2_xnor2_1 _2201_ (.Y(_0503_),
    .A(_0501_),
    .B(_0502_));
 sg13g2_xor2_1 _2202_ (.B(\u_usb_cdc.u_sie.data_q[3] ),
    .A(net548),
    .X(_0504_));
 sg13g2_xor2_1 _2203_ (.B(net762),
    .A(net563),
    .X(_0505_));
 sg13g2_xnor2_1 _2204_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_nor2b_1 _2205_ (.A(_0503_),
    .B_N(_0506_),
    .Y(_0507_));
 sg13g2_xnor2_1 _2206_ (.Y(_0508_),
    .A(_0503_),
    .B(_0506_));
 sg13g2_xor2_1 _2207_ (.B(\u_usb_cdc.u_sie.data_q[4] ),
    .A(\u_usb_cdc.u_sie.crc16_q[11] ),
    .X(_0509_));
 sg13g2_xor2_1 _2208_ (.B(net766),
    .A(net915),
    .X(_0510_));
 sg13g2_xnor2_1 _2209_ (.Y(_0511_),
    .A(\u_usb_cdc.u_sie.crc16_q[14] ),
    .B(net764));
 sg13g2_xnor2_1 _2210_ (.Y(_0512_),
    .A(_0510_),
    .B(_0511_));
 sg13g2_xnor2_1 _2211_ (.Y(_0513_),
    .A(_0509_),
    .B(_0512_));
 sg13g2_xnor2_1 _2212_ (.Y(_0514_),
    .A(_0508_),
    .B(_0513_));
 sg13g2_xnor2_1 _2213_ (.Y(_0515_),
    .A(_1946_),
    .B(_0512_));
 sg13g2_inv_1 _2214_ (.Y(_0516_),
    .A(_0515_));
 sg13g2_xnor2_1 _2215_ (.Y(_0517_),
    .A(net918),
    .B(_0510_));
 sg13g2_xnor2_1 _2216_ (.Y(_0518_),
    .A(_0504_),
    .B(_0509_));
 sg13g2_nand2_1 _2217_ (.Y(_0519_),
    .A(_0517_),
    .B(_0518_));
 sg13g2_xnor2_1 _2218_ (.Y(_0520_),
    .A(_0500_),
    .B(net541));
 sg13g2_xor2_1 _2219_ (.B(_0511_),
    .A(_0505_),
    .X(_0521_));
 sg13g2_inv_1 _2220_ (.Y(_0522_),
    .A(_0521_));
 sg13g2_xnor2_1 _2221_ (.Y(_0523_),
    .A(_0502_),
    .B(_0509_));
 sg13g2_nand4_1 _2222_ (.B(_1951_),
    .C(_1952_),
    .A(_1950_),
    .Y(_0524_),
    .D(_1953_));
 sg13g2_nor3_1 _2223_ (.A(\u_usb_cdc.u_sie.crc16_q[3] ),
    .B(\u_usb_cdc.u_sie.crc16_q[2] ),
    .C(_0524_),
    .Y(_0525_));
 sg13g2_nand3_1 _2224_ (.B(_0523_),
    .C(_0525_),
    .A(_0507_),
    .Y(_0526_));
 sg13g2_nor4_1 _2225_ (.A(_0519_),
    .B(_0520_),
    .C(_0522_),
    .D(_0526_),
    .Y(_0527_));
 sg13g2_and4_1 _2226_ (.A(_0500_),
    .B(_0514_),
    .C(_0516_),
    .D(_0527_),
    .X(_0528_));
 sg13g2_nand2_1 _2227_ (.Y(_0529_),
    .A(net706),
    .B(_0528_));
 sg13g2_a21oi_1 _2228_ (.A1(net833),
    .A2(_0529_),
    .Y(_0530_),
    .B1(net836));
 sg13g2_a21oi_1 _2229_ (.A1(_0499_),
    .A2(_0530_),
    .Y(_0531_),
    .B1(net746));
 sg13g2_xor2_1 _2230_ (.B(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .X(_0532_));
 sg13g2_xor2_1 _2231_ (.B(net779),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .X(_0533_));
 sg13g2_xor2_1 _2232_ (.B(net785),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .X(_0534_));
 sg13g2_xor2_1 _2233_ (.B(\u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .A(net775),
    .X(_0535_));
 sg13g2_xor2_1 _2234_ (.B(net772),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .X(_0536_));
 sg13g2_xor2_1 _2235_ (.B(net784),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .X(_0537_));
 sg13g2_xor2_1 _2236_ (.B(net787),
    .A(\u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .X(_0538_));
 sg13g2_nor3_1 _2237_ (.A(_0532_),
    .B(_0533_),
    .C(_0535_),
    .Y(_0539_));
 sg13g2_nor4_1 _2238_ (.A(_0534_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0540_));
 sg13g2_nand2b_2 _2239_ (.Y(_0541_),
    .B(net785),
    .A_N(net780));
 sg13g2_nand2b_2 _2240_ (.Y(_0542_),
    .B(_1915_),
    .A_N(_0541_));
 sg13g2_nor3_1 _2241_ (.A(net786),
    .B(net782),
    .C(net779),
    .Y(_0543_));
 sg13g2_nor2b_2 _2242_ (.A(net770),
    .B_N(net773),
    .Y(_0544_));
 sg13g2_nor2b_1 _2243_ (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .B_N(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .Y(_0545_));
 sg13g2_and4_1 _2244_ (.A(net785),
    .B(_0543_),
    .C(_0544_),
    .D(_0545_),
    .X(_0546_));
 sg13g2_nand2b_2 _2245_ (.Y(_0547_),
    .B(net787),
    .A_N(net782));
 sg13g2_nor2_2 _2246_ (.A(_1915_),
    .B(net715),
    .Y(_0548_));
 sg13g2_nand2_2 _2247_ (.Y(_0549_),
    .A(net786),
    .B(net785));
 sg13g2_nor2_2 _2248_ (.A(net781),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_nor3_2 _2249_ (.A(net780),
    .B(net777),
    .C(_0549_),
    .Y(_0551_));
 sg13g2_nor2_2 _2250_ (.A(net773),
    .B(net770),
    .Y(_0552_));
 sg13g2_and3_1 _2251_ (.X(_0553_),
    .A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .C(_0552_));
 sg13g2_a221oi_1 _2252_ (.B2(_0553_),
    .C1(_0546_),
    .B1(_0551_),
    .A1(_0539_),
    .Y(_0554_),
    .A2(_0540_));
 sg13g2_nor2b_1 _2253_ (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .B_N(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .Y(_0555_));
 sg13g2_nand2b_1 _2254_ (.Y(_0556_),
    .B(_0049_),
    .A_N(\u_usb_cdc.u_ctrl_endp.state_q[7] ));
 sg13g2_or4_1 _2255_ (.A(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .B(\u_usb_cdc.ctrl_stall ),
    .C(\u_usb_cdc.u_ctrl_endp.state_q[5] ),
    .D(_0556_),
    .X(_0557_));
 sg13g2_inv_1 _2256_ (.Y(_0558_),
    .A(_0557_));
 sg13g2_or2_1 _2257_ (.X(_0559_),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[1] ));
 sg13g2_nor3_1 _2258_ (.A(net841),
    .B(_0557_),
    .C(_0559_),
    .Y(_0560_));
 sg13g2_nor4_1 _2259_ (.A(net841),
    .B(_0555_),
    .C(_0557_),
    .D(_0559_),
    .Y(_0561_));
 sg13g2_or2_1 _2260_ (.X(_0562_),
    .B(net841),
    .A(net767));
 sg13g2_a21oi_1 _2261_ (.A1(_0554_),
    .A2(_0561_),
    .Y(_0563_),
    .B1(_0562_));
 sg13g2_nand2b_1 _2262_ (.Y(_0564_),
    .B(net803),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ));
 sg13g2_xnor2_1 _2263_ (.Y(_0565_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ),
    .B(net790));
 sg13g2_xnor2_1 _2264_ (.Y(_0566_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ),
    .B(net794));
 sg13g2_a22oi_1 _2265_ (.Y(_0567_),
    .B1(_1914_),
    .B2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ),
    .A2(_1912_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ));
 sg13g2_o21ai_1 _2266_ (.B1(_0567_),
    .Y(_0568_),
    .A1(_1914_),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ));
 sg13g2_nand4_1 _2267_ (.B(_0564_),
    .C(_0565_),
    .A(net767),
    .Y(_0569_),
    .D(_0566_));
 sg13g2_o21ai_1 _2268_ (.B1(net706),
    .Y(_0570_),
    .A1(_0568_),
    .A2(_0569_));
 sg13g2_nor2_1 _2269_ (.A(_0563_),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_and2_1 _2270_ (.A(_1906_),
    .B(net706),
    .X(_0572_));
 sg13g2_nand2_2 _2271_ (.Y(_0573_),
    .A(_1906_),
    .B(_1986_));
 sg13g2_nor2_1 _2272_ (.A(_1906_),
    .B(_1985_),
    .Y(_0574_));
 sg13g2_and2_1 _2273_ (.A(net767),
    .B(net706),
    .X(_0575_));
 sg13g2_nand2_2 _2274_ (.Y(_0576_),
    .A(net767),
    .B(net706));
 sg13g2_a221oi_1 _2275_ (.B2(net85),
    .C1(_0571_),
    .B1(net633),
    .A1(net165),
    .Y(_0577_),
    .A2(net634));
 sg13g2_nand2_2 _2276_ (.Y(_0578_),
    .A(net946),
    .B(net634));
 sg13g2_nand2b_2 _2277_ (.Y(_0579_),
    .B(_0578_),
    .A_N(_0577_));
 sg13g2_nand2_1 _2278_ (.Y(_0580_),
    .A(net839),
    .B(_0579_));
 sg13g2_and2_1 _2279_ (.A(net840),
    .B(_1989_),
    .X(_0581_));
 sg13g2_nor3_1 _2280_ (.A(\u_usb_cdc.u_sie.phy_state_q[2] ),
    .B(net186),
    .C(\u_usb_cdc.u_sie.phy_state_q[3] ),
    .Y(_0582_));
 sg13g2_a21oi_1 _2281_ (.A1(net208),
    .A2(_0582_),
    .Y(_0583_),
    .B1(net746));
 sg13g2_nor4_1 _2282_ (.A(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .B(net259),
    .C(_0581_),
    .D(_0583_),
    .Y(_0584_));
 sg13g2_nand2_2 _2283_ (.Y(_0585_),
    .A(_1993_),
    .B(net705));
 sg13g2_nand2b_1 _2284_ (.Y(_0586_),
    .B(_0053_),
    .A_N(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ));
 sg13g2_nand2b_1 _2285_ (.Y(_0587_),
    .B(_1997_),
    .A_N(_0586_));
 sg13g2_nor2_1 _2286_ (.A(_0585_),
    .B(_0587_),
    .Y(_0588_));
 sg13g2_nor3_2 _2287_ (.A(net746),
    .B(net748),
    .C(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq ),
    .Y(_0589_));
 sg13g2_o21ai_1 _2288_ (.B1(_0589_),
    .Y(_0590_),
    .A1(_0585_),
    .A2(_0587_));
 sg13g2_nand2_1 _2289_ (.Y(_0591_),
    .A(_1904_),
    .B(net743));
 sg13g2_and2_1 _2290_ (.A(net739),
    .B(_0590_),
    .X(_0592_));
 sg13g2_nand2_1 _2291_ (.Y(_0593_),
    .A(net743),
    .B(_0590_));
 sg13g2_nor2_1 _2292_ (.A(net747),
    .B(net596),
    .Y(_0594_));
 sg13g2_nand2_2 _2293_ (.Y(_0595_),
    .A(_1904_),
    .B(net597));
 sg13g2_nand3_1 _2294_ (.B(net260),
    .C(net592),
    .A(_0580_),
    .Y(_0596_));
 sg13g2_nand2_1 _2295_ (.Y(_0597_),
    .A(net208),
    .B(net595));
 sg13g2_nor2_1 _2296_ (.A(net746),
    .B(_0595_),
    .Y(_0598_));
 sg13g2_nor2_1 _2297_ (.A(_1903_),
    .B(_0528_),
    .Y(_0599_));
 sg13g2_nand2_1 _2298_ (.Y(_0600_),
    .A(net832),
    .B(net590));
 sg13g2_nor2b_2 _2299_ (.A(net745),
    .B_N(\u_usb_cdc.u_sie.phy_state_q[9] ),
    .Y(_0601_));
 sg13g2_nand4_1 _2300_ (.B(_0497_),
    .C(net591),
    .A(_0494_),
    .Y(_0602_),
    .D(_0601_));
 sg13g2_o21ai_1 _2301_ (.B1(_0597_),
    .Y(_0063_),
    .A1(_0531_),
    .A2(net261));
 sg13g2_nand2_1 _2302_ (.Y(_0603_),
    .A(net745),
    .B(_1904_));
 sg13g2_nand2_2 _2303_ (.Y(_0604_),
    .A(net745),
    .B(net833));
 sg13g2_nor2_2 _2304_ (.A(net747),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_nor2_2 _2305_ (.A(net749),
    .B(_0605_),
    .Y(_0606_));
 sg13g2_or2_1 _2306_ (.X(_0607_),
    .B(net749),
    .A(\u_usb_cdc.u_sie.out_eop_q ));
 sg13g2_nand4_1 _2307_ (.B(\u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .C(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .A(\u_usb_cdc.u_sie.delay_cnt_q[2] ),
    .Y(_0608_),
    .D(_0607_));
 sg13g2_nand2b_1 _2308_ (.Y(_0609_),
    .B(_0608_),
    .A_N(_0605_));
 sg13g2_and2_1 _2309_ (.A(net634),
    .B(_0609_),
    .X(_0610_));
 sg13g2_nand3_1 _2310_ (.B(net289),
    .C(net230),
    .A(net319),
    .Y(_0611_));
 sg13g2_nor3_1 _2311_ (.A(\u_usb_cdc.u_sie.in_byte_q[3] ),
    .B(_1989_),
    .C(_0611_),
    .Y(_0612_));
 sg13g2_nor4_1 _2312_ (.A(_1910_),
    .B(_0563_),
    .C(_0570_),
    .D(_0612_),
    .Y(_0613_));
 sg13g2_or3_1 _2313_ (.A(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .C(_0557_),
    .X(_0614_));
 sg13g2_nor2_1 _2314_ (.A(_0573_),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_nand2b_1 _2315_ (.Y(_0616_),
    .B(_0571_),
    .A_N(_0615_));
 sg13g2_inv_1 _2316_ (.Y(_0617_),
    .A(_0616_));
 sg13g2_nand2_1 _2317_ (.Y(_0618_),
    .A(net839),
    .B(_0578_));
 sg13g2_nor4_1 _2318_ (.A(_0563_),
    .B(_0570_),
    .C(_0615_),
    .D(_0618_),
    .Y(_0619_));
 sg13g2_o21ai_1 _2319_ (.B1(_0588_),
    .Y(_0620_),
    .A1(_0613_),
    .A2(_0619_));
 sg13g2_nor2_2 _2320_ (.A(\u_usb_cdc.sie_in_data_ack ),
    .B(\u_usb_cdc.sie_in_req ),
    .Y(_0621_));
 sg13g2_a21oi_1 _2321_ (.A1(_0620_),
    .A2(_0621_),
    .Y(_0622_),
    .B1(_0573_));
 sg13g2_nor2_2 _2322_ (.A(_1924_),
    .B(_0468_),
    .Y(_0623_));
 sg13g2_nand2_1 _2323_ (.Y(_0624_),
    .A(_0610_),
    .B(_0623_));
 sg13g2_o21ai_1 _2324_ (.B1(_0610_),
    .Y(_0625_),
    .A1(net749),
    .A2(_0623_));
 sg13g2_inv_1 _2325_ (.Y(_0626_),
    .A(_0625_));
 sg13g2_o21ai_1 _2326_ (.B1(_0625_),
    .Y(_0627_),
    .A1(_0610_),
    .A2(_0622_));
 sg13g2_nand2_1 _2327_ (.Y(_0628_),
    .A(\u_usb_cdc.sie_in_req ),
    .B(net634));
 sg13g2_o21ai_1 _2328_ (.B1(_0628_),
    .Y(_0629_),
    .A1(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .A2(\u_usb_cdc.u_ctrl_endp.state_q[5] ));
 sg13g2_a21oi_1 _2329_ (.A1(_1909_),
    .A2(net841),
    .Y(_0630_),
    .B1(\u_usb_cdc.u_ctrl_endp.state_q[2] ));
 sg13g2_a221oi_1 _2330_ (.B2(_0630_),
    .C1(_0573_),
    .B1(_0629_),
    .A1(_0620_),
    .Y(_0631_),
    .A2(_0621_));
 sg13g2_nor3_1 _2331_ (.A(net841),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[5] ),
    .C(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .Y(_0632_));
 sg13g2_nand2_1 _2332_ (.Y(_0633_),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .B(_0605_));
 sg13g2_nand2_1 _2333_ (.Y(_0634_),
    .A(_0632_),
    .B(_0633_));
 sg13g2_nand2_1 _2334_ (.Y(_0635_),
    .A(_0610_),
    .B(_0634_));
 sg13g2_nand2b_1 _2335_ (.Y(_0636_),
    .B(_0635_),
    .A_N(_0631_));
 sg13g2_nand3b_1 _2336_ (.B(_0635_),
    .C(net738),
    .Y(_0637_),
    .A_N(_0631_));
 sg13g2_nor2_2 _2337_ (.A(net588),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_or2_1 _2338_ (.X(_0639_),
    .B(net583),
    .A(net588));
 sg13g2_a21oi_1 _2339_ (.A1(\u_usb_cdc.sie_in_req ),
    .A2(net634),
    .Y(_0640_),
    .B1(\u_usb_cdc.sie_in_data_ack ));
 sg13g2_nand2_1 _2340_ (.Y(_0641_),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .B(_0640_));
 sg13g2_nand3b_1 _2341_ (.B(net535),
    .C(_0641_),
    .Y(_0642_),
    .A_N(\u_usb_cdc.u_ctrl_endp.state_q[3] ));
 sg13g2_nor2_1 _2342_ (.A(_0556_),
    .B(_0559_),
    .Y(_0643_));
 sg13g2_a21oi_1 _2343_ (.A1(_0632_),
    .A2(_0643_),
    .Y(_0644_),
    .B1(net714));
 sg13g2_nand3_1 _2344_ (.B(_0610_),
    .C(_0644_),
    .A(net750),
    .Y(_0645_));
 sg13g2_o21ai_1 _2345_ (.B1(net738),
    .Y(_0646_),
    .A1(_0610_),
    .A2(_0622_));
 sg13g2_inv_2 _2346_ (.Y(_0647_),
    .A(_0646_));
 sg13g2_o21ai_1 _2347_ (.B1(_0645_),
    .Y(_0648_),
    .A1(net535),
    .A2(_0647_));
 sg13g2_a21oi_1 _2348_ (.A1(_0638_),
    .A2(net536),
    .Y(_0062_),
    .B1(_0648_));
 sg13g2_nand2_2 _2349_ (.Y(_0649_),
    .A(_1917_),
    .B(_0552_));
 sg13g2_nor2b_2 _2350_ (.A(net777),
    .B_N(net782),
    .Y(_0650_));
 sg13g2_nand2_1 _2351_ (.Y(_0651_),
    .A(net786),
    .B(net715));
 sg13g2_nand3_1 _2352_ (.B(net715),
    .C(_0650_),
    .A(net786),
    .Y(_0652_));
 sg13g2_nor2_2 _2353_ (.A(net779),
    .B(_0649_),
    .Y(_0653_));
 sg13g2_or2_1 _2354_ (.X(_0654_),
    .B(_0649_),
    .A(net779));
 sg13g2_nand2_2 _2355_ (.Y(_0655_),
    .A(net784),
    .B(_0653_));
 sg13g2_inv_2 _2356_ (.Y(_0656_),
    .A(_0655_));
 sg13g2_nor2_1 _2357_ (.A(_0649_),
    .B(_0652_),
    .Y(_0657_));
 sg13g2_nand2_1 _2358_ (.Y(_0658_),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .B(_0605_));
 sg13g2_nor3_1 _2359_ (.A(net586),
    .B(net583),
    .C(net620),
    .Y(_0659_));
 sg13g2_nor2_1 _2360_ (.A(net786),
    .B(net785),
    .Y(_0660_));
 sg13g2_nand2_2 _2361_ (.Y(_0661_),
    .A(_1915_),
    .B(net716));
 sg13g2_nor2_2 _2362_ (.A(_0655_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_nand3_1 _2363_ (.B(_0656_),
    .C(_0659_),
    .A(net715),
    .Y(_0663_));
 sg13g2_nand2_1 _2364_ (.Y(_0664_),
    .A(net786),
    .B(net780));
 sg13g2_a21o_2 _2365_ (.A2(_0548_),
    .A1(net783),
    .B1(net778),
    .X(_0665_));
 sg13g2_nor2_1 _2366_ (.A(net773),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_nand4_1 _2367_ (.B(net785),
    .C(net783),
    .A(_1915_),
    .Y(_0667_),
    .D(net778));
 sg13g2_and2_1 _2368_ (.A(net774),
    .B(_0667_),
    .X(_0668_));
 sg13g2_nor2b_1 _2369_ (.A(net770),
    .B_N(net777),
    .Y(_0669_));
 sg13g2_nand2b_2 _2370_ (.Y(_0670_),
    .B(net776),
    .A_N(net774));
 sg13g2_nor2_1 _2371_ (.A(_0550_),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_nor4_1 _2372_ (.A(_0666_),
    .B(_0668_),
    .C(_0669_),
    .D(_0671_),
    .Y(_0672_));
 sg13g2_nand2b_2 _2373_ (.Y(_0673_),
    .B(_0672_),
    .A_N(_0649_));
 sg13g2_inv_1 _2374_ (.Y(_0674_),
    .A(_0673_));
 sg13g2_nor3_2 _2375_ (.A(net787),
    .B(net715),
    .C(_0655_),
    .Y(_0675_));
 sg13g2_nand2_1 _2376_ (.Y(_0676_),
    .A(net736),
    .B(_0675_));
 sg13g2_nor4_1 _2377_ (.A(net586),
    .B(net584),
    .C(net620),
    .D(_0676_),
    .Y(_0677_));
 sg13g2_a21oi_1 _2378_ (.A1(_0659_),
    .A2(_0674_),
    .Y(_0678_),
    .B1(_0677_));
 sg13g2_nor4_1 _2379_ (.A(net586),
    .B(net583),
    .C(_0653_),
    .D(net619),
    .Y(_0679_));
 sg13g2_or2_1 _2380_ (.X(_0680_),
    .B(net588),
    .A(net714));
 sg13g2_nor2b_2 _2381_ (.A(_0605_),
    .B_N(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .Y(_0681_));
 sg13g2_or4_1 _2382_ (.A(net841),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .C(_0557_),
    .D(_0681_),
    .X(_0682_));
 sg13g2_nor2_1 _2383_ (.A(net585),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_or4_1 _2384_ (.A(net714),
    .B(net588),
    .C(net585),
    .D(_0682_),
    .X(_0684_));
 sg13g2_nand2_1 _2385_ (.Y(_0685_),
    .A(_0550_),
    .B(_0653_));
 sg13g2_nand3_1 _2386_ (.B(_0550_),
    .C(_0653_),
    .A(net736),
    .Y(_0686_));
 sg13g2_nor4_1 _2387_ (.A(net586),
    .B(net584),
    .C(net619),
    .D(_0686_),
    .Y(_0687_));
 sg13g2_nor2_2 _2388_ (.A(_0542_),
    .B(_0654_),
    .Y(_0688_));
 sg13g2_inv_1 _2389_ (.Y(_0689_),
    .A(_0688_));
 sg13g2_nor4_1 _2390_ (.A(net587),
    .B(net583),
    .C(net619),
    .D(_0689_),
    .Y(_0690_));
 sg13g2_nor4_1 _2391_ (.A(_0679_),
    .B(_0684_),
    .C(_0687_),
    .D(_0690_),
    .Y(_0691_));
 sg13g2_nand3_1 _2392_ (.B(_0678_),
    .C(_0691_),
    .A(_0663_),
    .Y(_0692_));
 sg13g2_nor3_2 _2393_ (.A(net586),
    .B(net583),
    .C(net619),
    .Y(_0693_));
 sg13g2_nor4_1 _2394_ (.A(net586),
    .B(net583),
    .C(net620),
    .D(_0673_),
    .Y(_0694_));
 sg13g2_nor3_2 _2395_ (.A(net587),
    .B(net584),
    .C(net620),
    .Y(_0695_));
 sg13g2_nor4_1 _2396_ (.A(net586),
    .B(net584),
    .C(net619),
    .D(_0686_),
    .Y(_0696_));
 sg13g2_nand2_1 _2397_ (.Y(_0697_),
    .A(net738),
    .B(_0688_));
 sg13g2_nor4_2 _2398_ (.A(net587),
    .B(net584),
    .C(net619),
    .Y(_0698_),
    .D(_0697_));
 sg13g2_nand2_1 _2399_ (.Y(_0699_),
    .A(_0675_),
    .B(net574));
 sg13g2_nand2_1 _2400_ (.Y(_0700_),
    .A(_0662_),
    .B(net574));
 sg13g2_or4_1 _2401_ (.A(net841),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .C(_0557_),
    .D(_0681_),
    .X(_0701_));
 sg13g2_nor2_2 _2402_ (.A(net755),
    .B(\u_usb_cdc.sie_out_data[2] ),
    .Y(_0702_));
 sg13g2_nand2_1 _2403_ (.Y(_0703_),
    .A(_0478_),
    .B(_0702_));
 sg13g2_nand4_1 _2404_ (.B(_1901_),
    .C(_0478_),
    .A(_1899_),
    .Y(_0704_),
    .D(_0702_));
 sg13g2_nor2_2 _2405_ (.A(net784),
    .B(_0661_),
    .Y(_0705_));
 sg13g2_nor4_1 _2406_ (.A(net784),
    .B(_0654_),
    .C(_0661_),
    .D(_0704_),
    .Y(_0706_));
 sg13g2_a22oi_1 _2407_ (.Y(_0061_),
    .B1(net574),
    .B2(_0706_),
    .A2(_0692_),
    .A1(_1982_));
 sg13g2_and2_1 _2408_ (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .B(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .X(\u_usb_cdc.configured_o ));
 sg13g2_nor4_2 _2409_ (.A(net753),
    .B(net754),
    .C(net751),
    .Y(_0707_),
    .D(net752));
 sg13g2_nand2_1 _2410_ (.Y(_0708_),
    .A(_0702_),
    .B(_0707_));
 sg13g2_nor2_1 _2411_ (.A(net757),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_nand3_1 _2412_ (.B(_0702_),
    .C(_0707_),
    .A(net720),
    .Y(_0710_));
 sg13g2_nor2_1 _2413_ (.A(net760),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_nand4_1 _2414_ (.B(_0656_),
    .C(_0659_),
    .A(net715),
    .Y(_0712_),
    .D(net617));
 sg13g2_nor2_2 _2415_ (.A(net721),
    .B(_0710_),
    .Y(_0713_));
 sg13g2_nand2_1 _2416_ (.Y(_0714_),
    .A(net760),
    .B(_0709_));
 sg13g2_nand3_1 _2417_ (.B(_0656_),
    .C(net574),
    .A(net715),
    .Y(_0715_));
 sg13g2_nand4_1 _2418_ (.B(_0656_),
    .C(net574),
    .A(net715),
    .Y(_0716_),
    .D(net617));
 sg13g2_or4_1 _2419_ (.A(net714),
    .B(net586),
    .C(net584),
    .D(_0701_),
    .X(_0717_));
 sg13g2_a221oi_1 _2420_ (.B2(net617),
    .C1(_0717_),
    .B1(_0698_),
    .A1(_0654_),
    .Y(_0718_),
    .A2(net574));
 sg13g2_o21ai_1 _2421_ (.B1(net617),
    .Y(_0719_),
    .A1(_0694_),
    .A2(_0696_));
 sg13g2_nand3_1 _2422_ (.B(_0718_),
    .C(_0719_),
    .A(_0716_),
    .Y(_0720_));
 sg13g2_nor2_1 _2423_ (.A(_0699_),
    .B(_0714_),
    .Y(_0721_));
 sg13g2_nand3_1 _2424_ (.B(_0693_),
    .C(_0713_),
    .A(_0675_),
    .Y(_0722_));
 sg13g2_nor3_1 _2425_ (.A(net588),
    .B(net585),
    .C(_0682_),
    .Y(_0723_));
 sg13g2_nand2_2 _2426_ (.Y(_0724_),
    .A(net738),
    .B(_0723_));
 sg13g2_o21ai_1 _2427_ (.B1(net971),
    .Y(_0725_),
    .A1(_0720_),
    .A2(_0721_));
 sg13g2_nand2b_2 _2428_ (.Y(_0726_),
    .B(net937),
    .A_N(net346));
 sg13g2_nand2_1 _2429_ (.Y(_0727_),
    .A(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .B(_0726_));
 sg13g2_nand3_1 _2430_ (.B(_1927_),
    .C(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .A(_1926_),
    .Y(_0728_));
 sg13g2_nor2b_1 _2431_ (.A(_0728_),
    .B_N(_0726_),
    .Y(_0729_));
 sg13g2_nand3_1 _2432_ (.B(net718),
    .C(_0707_),
    .A(net1016),
    .Y(_0730_));
 sg13g2_nor3_1 _2433_ (.A(net760),
    .B(net757),
    .C(_0730_),
    .Y(_0731_));
 sg13g2_nand2_1 _2434_ (.Y(_0732_),
    .A(_0729_),
    .B(_0731_));
 sg13g2_nand2_1 _2435_ (.Y(_0733_),
    .A(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .B(_0624_));
 sg13g2_or2_1 _2436_ (.X(_0734_),
    .B(_0733_),
    .A(net584));
 sg13g2_nor3_2 _2437_ (.A(net747),
    .B(net750),
    .C(_0604_),
    .Y(_0735_));
 sg13g2_nand2_2 _2438_ (.Y(_0736_),
    .A(net634),
    .B(_0735_));
 sg13g2_or3_1 _2439_ (.A(net884),
    .B(_0734_),
    .C(_0736_),
    .X(_0737_));
 sg13g2_nor2_1 _2440_ (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .B(_0547_),
    .Y(_0738_));
 sg13g2_nand3_1 _2441_ (.B(_0653_),
    .C(_0738_),
    .A(net736),
    .Y(_0739_));
 sg13g2_nor2_1 _2442_ (.A(net860),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_nand2b_2 _2443_ (.Y(_0741_),
    .B(_0740_),
    .A_N(_0737_));
 sg13g2_o21ai_1 _2444_ (.B1(_0725_),
    .Y(_0005_),
    .A1(_0732_),
    .A2(_0741_));
 sg13g2_nand2_1 _2445_ (.Y(_0742_),
    .A(net953),
    .B(_0692_));
 sg13g2_nor2_2 _2446_ (.A(_0480_),
    .B(_0708_),
    .Y(_0743_));
 sg13g2_nor4_1 _2447_ (.A(net755),
    .B(net756),
    .C(\u_usb_cdc.sie_out_data[4] ),
    .D(net752),
    .Y(_0744_));
 sg13g2_and4_1 _2448_ (.A(\u_usb_cdc.sie_out_data[5] ),
    .B(net717),
    .C(\u_usb_cdc.configured_o ),
    .D(_0744_),
    .X(_0745_));
 sg13g2_nor2_1 _2449_ (.A(_0739_),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_or2_1 _2450_ (.X(_0747_),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[4] ));
 sg13g2_nor2_1 _2451_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .B(net842),
    .Y(_0748_));
 sg13g2_nor3_1 _2452_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .B(net842),
    .C(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .Y(_0749_));
 sg13g2_inv_1 _2453_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_nor3_1 _2454_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .B(_0747_),
    .C(_0750_),
    .Y(_0751_));
 sg13g2_nor2_2 _2455_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .Y(_0752_));
 sg13g2_nor3_1 _2456_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .B(net842),
    .C(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .Y(_0753_));
 sg13g2_nand2_1 _2457_ (.Y(_0754_),
    .A(_0752_),
    .B(_0753_));
 sg13g2_nor3_1 _2458_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .C(_0747_),
    .Y(_0755_));
 sg13g2_inv_1 _2459_ (.Y(_0756_),
    .A(_0755_));
 sg13g2_a21oi_1 _2460_ (.A1(_0673_),
    .A2(_0685_),
    .Y(_0757_),
    .B1(_0751_));
 sg13g2_nand2_1 _2461_ (.Y(_0758_),
    .A(_0751_),
    .B(_0752_));
 sg13g2_a22oi_1 _2462_ (.Y(_0759_),
    .B1(_0758_),
    .B2(_0657_),
    .A2(_0756_),
    .A1(_0688_));
 sg13g2_a21oi_1 _2463_ (.A1(_0662_),
    .A2(_0754_),
    .Y(_0760_),
    .B1(_0757_));
 sg13g2_a21oi_1 _2464_ (.A1(_0759_),
    .A2(_0760_),
    .Y(_0761_),
    .B1(net617));
 sg13g2_nand3_1 _2465_ (.B(_0714_),
    .C(_0747_),
    .A(_0675_),
    .Y(_0762_));
 sg13g2_nand3_1 _2466_ (.B(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .C(net618),
    .A(_1926_),
    .Y(_0763_));
 sg13g2_nand3_1 _2467_ (.B(_0688_),
    .C(_0763_),
    .A(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .Y(_0764_));
 sg13g2_nand3_1 _2468_ (.B(_0704_),
    .C(_0705_),
    .A(_0653_),
    .Y(_0765_));
 sg13g2_nor2_1 _2469_ (.A(net720),
    .B(net751),
    .Y(_0766_));
 sg13g2_nor4_1 _2470_ (.A(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .B(_1927_),
    .C(_0703_),
    .D(_0766_),
    .Y(_0767_));
 sg13g2_a21oi_1 _2471_ (.A1(net760),
    .A2(_1926_),
    .Y(_0768_),
    .B1(_0710_));
 sg13g2_a21oi_1 _2472_ (.A1(_1927_),
    .A2(_0768_),
    .Y(_0769_),
    .B1(_0767_));
 sg13g2_a22oi_1 _2473_ (.Y(_0770_),
    .B1(_0769_),
    .B2(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .A2(_0710_),
    .A1(\u_usb_cdc.u_ctrl_endp.req_q[11] ));
 sg13g2_o21ai_1 _2474_ (.B1(_0770_),
    .Y(_0771_),
    .A1(_1931_),
    .A2(_0767_));
 sg13g2_nand2_1 _2475_ (.Y(_0772_),
    .A(_0662_),
    .B(_0771_));
 sg13g2_nand4_1 _2476_ (.B(_0764_),
    .C(_0765_),
    .A(_0762_),
    .Y(_0773_),
    .D(_0772_));
 sg13g2_o21ai_1 _2477_ (.B1(net736),
    .Y(_0774_),
    .A1(_0761_),
    .A2(_0773_));
 sg13g2_nor3_1 _2478_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .C(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .Y(_0775_));
 sg13g2_nand3_1 _2479_ (.B(_0752_),
    .C(_0775_),
    .A(_0751_),
    .Y(_0776_));
 sg13g2_nand2b_1 _2480_ (.Y(_0777_),
    .B(_0776_),
    .A_N(_0739_));
 sg13g2_nand3_1 _2481_ (.B(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .C(_0688_),
    .A(net738),
    .Y(_0778_));
 sg13g2_or2_1 _2482_ (.X(_0779_),
    .B(_0778_),
    .A(net717));
 sg13g2_nor2_1 _2483_ (.A(_1933_),
    .B(_0686_),
    .Y(_0780_));
 sg13g2_nor4_1 _2484_ (.A(_1933_),
    .B(_0686_),
    .C(_0713_),
    .D(_0743_),
    .Y(_0781_));
 sg13g2_nor2_1 _2485_ (.A(_0676_),
    .B(_0747_),
    .Y(_0782_));
 sg13g2_nor4_1 _2486_ (.A(_0676_),
    .B(net617),
    .C(_0747_),
    .D(_0749_),
    .Y(_0783_));
 sg13g2_nand3_1 _2487_ (.B(net842),
    .C(_0688_),
    .A(net738),
    .Y(_0784_));
 sg13g2_nor2_1 _2488_ (.A(_0709_),
    .B(_0784_),
    .Y(_0785_));
 sg13g2_nor3_1 _2489_ (.A(_0781_),
    .B(_0783_),
    .C(_0785_),
    .Y(_0786_));
 sg13g2_nand4_1 _2490_ (.B(_0777_),
    .C(_0779_),
    .A(_0774_),
    .Y(_0787_),
    .D(_0786_));
 sg13g2_nand3_1 _2491_ (.B(\u_usb_cdc.sie_out_data[2] ),
    .C(_0707_),
    .A(net719),
    .Y(_0788_));
 sg13g2_nor2_1 _2492_ (.A(_0480_),
    .B(_0788_),
    .Y(_0789_));
 sg13g2_a221oi_1 _2493_ (.B2(_0789_),
    .C1(_0731_),
    .B1(_0728_),
    .A1(net618),
    .Y(_0790_),
    .A2(_0727_));
 sg13g2_or2_1 _2494_ (.X(_0791_),
    .B(_0790_),
    .A(_0729_));
 sg13g2_o21ai_1 _2495_ (.B1(_0730_),
    .Y(_0792_),
    .A1(_0479_),
    .A2(_0788_));
 sg13g2_nor2_1 _2496_ (.A(_0709_),
    .B(_0792_),
    .Y(_0793_));
 sg13g2_nand4_1 _2497_ (.B(_1927_),
    .C(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .A(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .Y(_0794_),
    .D(\u_usb_cdc.configured_o ));
 sg13g2_nor2_1 _2498_ (.A(_0480_),
    .B(_0730_),
    .Y(_0795_));
 sg13g2_a221oi_1 _2499_ (.B2(_0795_),
    .C1(_0793_),
    .B1(_0794_),
    .A1(net760),
    .Y(_0796_),
    .A2(net758));
 sg13g2_a21oi_1 _2500_ (.A1(_0791_),
    .A2(_0796_),
    .Y(_0797_),
    .B1(_0739_));
 sg13g2_nor3_1 _2501_ (.A(net920),
    .B(net910),
    .C(net993),
    .Y(_0798_));
 sg13g2_inv_1 _2502_ (.Y(_0799_),
    .A(_0798_));
 sg13g2_nor3_1 _2503_ (.A(net721),
    .B(net757),
    .C(_0739_),
    .Y(_0800_));
 sg13g2_nand2b_1 _2504_ (.Y(_0801_),
    .B(_0800_),
    .A_N(_0788_));
 sg13g2_nand2b_1 _2505_ (.Y(_0802_),
    .B(_0800_),
    .A_N(_0730_));
 sg13g2_and2_1 _2506_ (.A(_1928_),
    .B(_0726_),
    .X(_0803_));
 sg13g2_nor3_1 _2507_ (.A(_0714_),
    .B(_0739_),
    .C(_0803_),
    .Y(_0804_));
 sg13g2_nor2_1 _2508_ (.A(_0726_),
    .B(_0802_),
    .Y(_0805_));
 sg13g2_a21oi_1 _2509_ (.A1(_0801_),
    .A2(_0802_),
    .Y(_0806_),
    .B1(_0798_));
 sg13g2_nor4_1 _2510_ (.A(_0797_),
    .B(_0804_),
    .C(_0805_),
    .D(_0806_),
    .Y(_0807_));
 sg13g2_nor4_1 _2511_ (.A(net884),
    .B(_0734_),
    .C(_0736_),
    .D(_0807_),
    .Y(_0808_));
 sg13g2_a21oi_1 _2512_ (.A1(_0695_),
    .A2(_0787_),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_nor3_1 _2513_ (.A(_1930_),
    .B(_0699_),
    .C(_0743_),
    .Y(_0810_));
 sg13g2_nor3_1 _2514_ (.A(_1905_),
    .B(_0734_),
    .C(_0736_),
    .Y(_0811_));
 sg13g2_a21oi_1 _2515_ (.A1(_0746_),
    .A2(_0811_),
    .Y(_0812_),
    .B1(_0810_));
 sg13g2_nand3_1 _2516_ (.B(_0809_),
    .C(_0812_),
    .A(_0742_),
    .Y(_0004_));
 sg13g2_nand2_1 _2517_ (.Y(_0813_),
    .A(_0698_),
    .B(_0713_));
 sg13g2_nand3_1 _2518_ (.B(net618),
    .C(_0782_),
    .A(_0695_),
    .Y(_0814_));
 sg13g2_nand2_1 _2519_ (.Y(_0815_),
    .A(_0813_),
    .B(_0814_));
 sg13g2_o21ai_1 _2520_ (.B1(net842),
    .Y(_0816_),
    .A1(_0720_),
    .A2(_0815_));
 sg13g2_nor4_1 _2521_ (.A(net884),
    .B(net860),
    .C(_0734_),
    .D(_0736_),
    .Y(_0817_));
 sg13g2_nand3_1 _2522_ (.B(_0798_),
    .C(_0817_),
    .A(_0726_),
    .Y(_0818_));
 sg13g2_o21ai_1 _2523_ (.B1(_0816_),
    .Y(_0006_),
    .A1(_0802_),
    .A2(_0818_));
 sg13g2_or2_1 _2524_ (.X(_0819_),
    .B(_0683_),
    .A(_0680_));
 sg13g2_nand3_1 _2525_ (.B(_0814_),
    .C(_0819_),
    .A(_0719_),
    .Y(_0820_));
 sg13g2_nor2_1 _2526_ (.A(_0679_),
    .B(_0680_),
    .Y(_0821_));
 sg13g2_nand4_1 _2527_ (.B(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .C(_0698_),
    .A(_1926_),
    .Y(_0822_),
    .D(net618));
 sg13g2_nand3_1 _2528_ (.B(net574),
    .C(net617),
    .A(_0657_),
    .Y(_0823_));
 sg13g2_nand3_1 _2529_ (.B(_0693_),
    .C(_0767_),
    .A(_0662_),
    .Y(_0824_));
 sg13g2_nand4_1 _2530_ (.B(_0822_),
    .C(_0823_),
    .A(_0821_),
    .Y(_0825_),
    .D(_0824_));
 sg13g2_o21ai_1 _2531_ (.B1(net906),
    .Y(_0826_),
    .A1(_0820_),
    .A2(_0825_));
 sg13g2_nand2_1 _2532_ (.Y(_0827_),
    .A(_0713_),
    .B(_0803_));
 sg13g2_o21ai_1 _2533_ (.B1(_0826_),
    .Y(_0007_),
    .A1(_0741_),
    .A2(_0827_));
 sg13g2_nand2_1 _2534_ (.Y(_0828_),
    .A(net717),
    .B(_0698_));
 sg13g2_nand3_1 _2535_ (.B(_0821_),
    .C(_0828_),
    .A(_0712_),
    .Y(_0829_));
 sg13g2_o21ai_1 _2536_ (.B1(net921),
    .Y(_0830_),
    .A1(_0820_),
    .A2(_0829_));
 sg13g2_or4_1 _2537_ (.A(net860),
    .B(_0737_),
    .C(_0799_),
    .D(_0801_),
    .X(_0831_));
 sg13g2_nand2_1 _2538_ (.Y(_0008_),
    .A(_0830_),
    .B(_0831_));
 sg13g2_nand3_1 _2539_ (.B(_0691_),
    .C(_0712_),
    .A(_0678_),
    .Y(_0832_));
 sg13g2_nand2_1 _2540_ (.Y(_0833_),
    .A(net845),
    .B(_0832_));
 sg13g2_nand3_1 _2541_ (.B(_0743_),
    .C(_0780_),
    .A(_0695_),
    .Y(_0834_));
 sg13g2_nand2_1 _2542_ (.Y(_0009_),
    .A(_0833_),
    .B(_0834_));
 sg13g2_o21ai_1 _2543_ (.B1(net574),
    .Y(_0835_),
    .A1(_0674_),
    .A2(_0675_));
 sg13g2_nand3_1 _2544_ (.B(_0718_),
    .C(_0835_),
    .A(_0715_),
    .Y(_0836_));
 sg13g2_nor4_1 _2545_ (.A(_0480_),
    .B(_0728_),
    .C(_0741_),
    .D(_0788_),
    .Y(_0837_));
 sg13g2_a21o_1 _2546_ (.A2(_0836_),
    .A1(net949),
    .B1(_0837_),
    .X(_0010_));
 sg13g2_nand2_1 _2547_ (.Y(_0838_),
    .A(net206),
    .B(_0692_));
 sg13g2_nand3_1 _2548_ (.B(_0745_),
    .C(_0811_),
    .A(_0740_),
    .Y(_0839_));
 sg13g2_nand2_1 _2549_ (.Y(_0000_),
    .A(_0838_),
    .B(_0839_));
 sg13g2_nand3_1 _2550_ (.B(_0719_),
    .C(_0823_),
    .A(_0718_),
    .Y(_0840_));
 sg13g2_o21ai_1 _2551_ (.B1(_0722_),
    .Y(_0841_),
    .A1(_0700_),
    .A2(_0710_));
 sg13g2_o21ai_1 _2552_ (.B1(net552),
    .Y(_0842_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_nand2b_1 _2553_ (.Y(_0843_),
    .B(_0795_),
    .A_N(_0794_));
 sg13g2_o21ai_1 _2554_ (.B1(_0842_),
    .Y(_0001_),
    .A1(_0741_),
    .A2(_0843_));
 sg13g2_or2_1 _2555_ (.X(_0844_),
    .B(net585),
    .A(_0626_));
 sg13g2_nor2b_1 _2556_ (.A(_0844_),
    .B_N(_0628_),
    .Y(_0845_));
 sg13g2_o21ai_1 _2557_ (.B1(net550),
    .Y(_0846_),
    .A1(_0646_),
    .A2(_0845_));
 sg13g2_or2_1 _2558_ (.X(_0847_),
    .B(net854),
    .A(net538));
 sg13g2_or4_1 _2559_ (.A(net864),
    .B(net856),
    .C(net523),
    .D(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .X(_0848_));
 sg13g2_nor3_1 _2560_ (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .B(_0847_),
    .C(_0848_),
    .Y(_0849_));
 sg13g2_nand2_1 _2561_ (.Y(_0850_),
    .A(net779),
    .B(_0705_));
 sg13g2_nor3_1 _2562_ (.A(net953),
    .B(_0649_),
    .C(_0850_),
    .Y(_0851_));
 sg13g2_inv_1 _2563_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_nand4_1 _2564_ (.B(_0638_),
    .C(_0681_),
    .A(_1928_),
    .Y(_0853_),
    .D(_0851_));
 sg13g2_o21ai_1 _2565_ (.B1(_0846_),
    .Y(_0011_),
    .A1(_0849_),
    .A2(_0853_));
 sg13g2_nor3_1 _2566_ (.A(net750),
    .B(_0624_),
    .C(_0646_),
    .Y(_0854_));
 sg13g2_a221oi_1 _2567_ (.B2(net739),
    .C1(_0854_),
    .B1(_0695_),
    .A1(net1037),
    .Y(_0855_),
    .A2(_0646_));
 sg13g2_inv_1 _2568_ (.Y(_0012_),
    .A(net1038));
 sg13g2_nor2_1 _2569_ (.A(_0626_),
    .B(_0628_),
    .Y(_0856_));
 sg13g2_nand2_1 _2570_ (.Y(_0857_),
    .A(net550),
    .B(_0856_));
 sg13g2_a22oi_1 _2571_ (.Y(_0858_),
    .B1(_0646_),
    .B2(net871),
    .A2(_0638_),
    .A1(net866));
 sg13g2_o21ai_1 _2572_ (.B1(_0858_),
    .Y(_0013_),
    .A1(net583),
    .A2(_0857_));
 sg13g2_nand2b_1 _2573_ (.Y(_0859_),
    .B(net946),
    .A_N(_0854_));
 sg13g2_a21oi_1 _2574_ (.A1(_0681_),
    .A2(_0852_),
    .Y(_0860_),
    .B1(net584));
 sg13g2_o21ai_1 _2575_ (.B1(net947),
    .Y(_0014_),
    .A1(_0680_),
    .A2(_0860_));
 sg13g2_or4_1 _2576_ (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .B(_0847_),
    .C(_0848_),
    .D(_0853_),
    .X(_0861_));
 sg13g2_o21ai_1 _2577_ (.B1(_0861_),
    .Y(_0015_),
    .A1(_1919_),
    .A2(_0647_));
 sg13g2_nor3_1 _2578_ (.A(\u_usb_cdc.sie_in_data_ack ),
    .B(_0554_),
    .C(net583),
    .Y(_0862_));
 sg13g2_a221oi_1 _2579_ (.B2(_0862_),
    .C1(_0646_),
    .B1(_0856_),
    .A1(_0554_),
    .Y(_0863_),
    .A2(_0638_));
 sg13g2_nand4_1 _2580_ (.B(_0638_),
    .C(_0681_),
    .A(net993),
    .Y(_0864_),
    .D(_0851_));
 sg13g2_o21ai_1 _2581_ (.B1(_0864_),
    .Y(_0016_),
    .A1(_1920_),
    .A2(_0863_));
 sg13g2_nor2_1 _2582_ (.A(_1920_),
    .B(_0554_),
    .Y(_0865_));
 sg13g2_a21oi_1 _2583_ (.A1(\u_usb_cdc.sie_in_data_ack ),
    .A2(_0865_),
    .Y(_0866_),
    .B1(net888));
 sg13g2_nor3_1 _2584_ (.A(_0639_),
    .B(_0640_),
    .C(_0866_),
    .Y(_0867_));
 sg13g2_a21o_1 _2585_ (.A2(_0646_),
    .A1(net888),
    .B1(_0867_),
    .X(_0017_));
 sg13g2_nand2_1 _2586_ (.Y(_0868_),
    .A(net840),
    .B(net595));
 sg13g2_nand4_1 _2587_ (.B(_0496_),
    .C(net590),
    .A(_0494_),
    .Y(_0869_),
    .D(_0601_));
 sg13g2_nor2_1 _2588_ (.A(net745),
    .B(_0498_),
    .Y(_0870_));
 sg13g2_o21ai_1 _2589_ (.B1(_0868_),
    .Y(_0020_),
    .A1(_0469_),
    .A2(net582));
 sg13g2_nand2_1 _2590_ (.Y(_0871_),
    .A(net413),
    .B(net595));
 sg13g2_nand2_1 _2591_ (.Y(_0872_),
    .A(net746),
    .B(net592));
 sg13g2_nand3_1 _2592_ (.B(net837),
    .C(net592),
    .A(net746),
    .Y(_0873_));
 sg13g2_xor2_1 _2593_ (.B(\u_usb_cdc.u_sie.addr_q[2] ),
    .A(\u_usb_cdc.addr[2] ),
    .X(_0874_));
 sg13g2_xnor2_1 _2594_ (.Y(_0875_),
    .A(\u_usb_cdc.addr[1] ),
    .B(net252));
 sg13g2_xor2_1 _2595_ (.B(\u_usb_cdc.u_sie.addr_q[5] ),
    .A(\u_usb_cdc.addr[5] ),
    .X(_0876_));
 sg13g2_xnor2_1 _2596_ (.Y(_0877_),
    .A(\u_usb_cdc.addr[3] ),
    .B(net200));
 sg13g2_xor2_1 _2597_ (.B(\u_usb_cdc.u_sie.addr_q[0] ),
    .A(\u_usb_cdc.addr[0] ),
    .X(_0878_));
 sg13g2_xnor2_1 _2598_ (.Y(_0879_),
    .A(\u_usb_cdc.addr[6] ),
    .B(net250));
 sg13g2_xor2_1 _2599_ (.B(\u_usb_cdc.u_sie.addr_q[4] ),
    .A(\u_usb_cdc.addr[4] ),
    .X(_0880_));
 sg13g2_nor4_1 _2600_ (.A(_0874_),
    .B(_0876_),
    .C(_0878_),
    .D(_0880_),
    .Y(_0881_));
 sg13g2_nand4_1 _2601_ (.B(_0877_),
    .C(_0879_),
    .A(_0875_),
    .Y(_0882_),
    .D(_0881_));
 sg13g2_a21oi_1 _2602_ (.A1(_1924_),
    .A2(\u_usb_cdc.u_sie.pid_q[3] ),
    .Y(_0883_),
    .B1(net762));
 sg13g2_nand4_1 _2603_ (.B(_0467_),
    .C(_0495_),
    .A(net706),
    .Y(_0884_),
    .D(_0883_));
 sg13g2_xnor2_1 _2604_ (.Y(_0885_),
    .A(net766),
    .B(\u_usb_cdc.u_sie.data_q[4] ));
 sg13g2_xnor2_1 _2605_ (.Y(_0886_),
    .A(net764),
    .B(\u_usb_cdc.u_sie.data_q[5] ));
 sg13g2_xnor2_1 _2606_ (.Y(_0887_),
    .A(\u_usb_cdc.u_sie.data_q[3] ),
    .B(\u_usb_cdc.u_sie.data_q[7] ));
 sg13g2_xnor2_1 _2607_ (.Y(_0888_),
    .A(net762),
    .B(\u_usb_cdc.u_sie.data_q[6] ));
 sg13g2_nor4_2 _2608_ (.A(_0885_),
    .B(_0886_),
    .C(_0887_),
    .Y(_0889_),
    .D(_0888_));
 sg13g2_nand2_2 _2609_ (.Y(_0890_),
    .A(net766),
    .B(_0889_));
 sg13g2_nor3_1 _2610_ (.A(_0882_),
    .B(_0884_),
    .C(_0890_),
    .Y(_0891_));
 sg13g2_nand2_1 _2611_ (.Y(_0892_),
    .A(net764),
    .B(_0891_));
 sg13g2_o21ai_1 _2612_ (.B1(_0871_),
    .Y(_0021_),
    .A1(_0873_),
    .A2(_0892_));
 sg13g2_nor3_1 _2613_ (.A(net764),
    .B(_0873_),
    .C(_0890_),
    .Y(_0893_));
 sg13g2_a21o_1 _2614_ (.A2(net595),
    .A1(net525),
    .B1(_0893_),
    .X(_0022_));
 sg13g2_nand2_2 _2615_ (.Y(_0894_),
    .A(net835),
    .B(net592));
 sg13g2_nand2_1 _2616_ (.Y(_0895_),
    .A(_1990_),
    .B(_0578_));
 sg13g2_or2_1 _2617_ (.X(_0896_),
    .B(_0895_),
    .A(_0595_));
 sg13g2_nor3_1 _2618_ (.A(_0577_),
    .B(_0617_),
    .C(_0896_),
    .Y(_0897_));
 sg13g2_a21oi_1 _2619_ (.A1(net838),
    .A2(net593),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_o21ai_1 _2620_ (.B1(_0898_),
    .Y(_0023_),
    .A1(_0613_),
    .A2(_0894_));
 sg13g2_o21ai_1 _2621_ (.B1(net837),
    .Y(_0899_),
    .A1(net764),
    .A2(_0890_));
 sg13g2_nor2_1 _2622_ (.A(_0891_),
    .B(_0899_),
    .Y(_0900_));
 sg13g2_o21ai_1 _2623_ (.B1(_0592_),
    .Y(_0901_),
    .A1(net832),
    .A2(_0900_));
 sg13g2_a22oi_1 _2624_ (.Y(_0024_),
    .B1(_0901_),
    .B2(_1956_),
    .A2(_0603_),
    .A1(_0592_));
 sg13g2_nand2_1 _2625_ (.Y(_0902_),
    .A(net837),
    .B(net595));
 sg13g2_o21ai_1 _2626_ (.B1(_0902_),
    .Y(_0025_),
    .A1(net208),
    .A2(_0872_));
 sg13g2_a22oi_1 _2627_ (.Y(_0903_),
    .B1(_0613_),
    .B2(_1904_),
    .A2(net593),
    .A1(net835));
 sg13g2_o21ai_1 _2628_ (.B1(_0903_),
    .Y(_0026_),
    .A1(_0616_),
    .A2(_0896_));
 sg13g2_nand2_1 _2629_ (.Y(_0904_),
    .A(net847),
    .B(net595));
 sg13g2_nor2_2 _2630_ (.A(net847),
    .B(net413),
    .Y(_0905_));
 sg13g2_o21ai_1 _2631_ (.B1(_0904_),
    .Y(_0027_),
    .A1(_0872_),
    .A2(_0905_));
 sg13g2_nand2_1 _2632_ (.Y(_0906_),
    .A(net832),
    .B(net595));
 sg13g2_o21ai_1 _2633_ (.B1(_0906_),
    .Y(_0028_),
    .A1(_1957_),
    .A2(_0872_));
 sg13g2_a22oi_1 _2634_ (.Y(_0907_),
    .B1(net592),
    .B2(net939),
    .A2(net596),
    .A1(net259));
 sg13g2_inv_1 _2635_ (.Y(_0018_),
    .A(_0907_));
 sg13g2_nor2_1 _2636_ (.A(net745),
    .B(_1903_),
    .Y(_0908_));
 sg13g2_nor2b_1 _2637_ (.A(_0529_),
    .B_N(_0908_),
    .Y(_0909_));
 sg13g2_a22oi_1 _2638_ (.Y(_0910_),
    .B1(net592),
    .B2(_0909_),
    .A2(net595),
    .A1(net975));
 sg13g2_inv_1 _2639_ (.Y(_0019_),
    .A(_0910_));
 sg13g2_nor2_1 _2640_ (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[2] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ),
    .Y(_0911_));
 sg13g2_nor4_1 _2641_ (.A(_0056_),
    .B(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .C(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ),
    .D(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .Y(_0912_));
 sg13g2_nand4_1 _2642_ (.B(_0446_),
    .C(_0911_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ),
    .Y(_0913_),
    .D(_0912_));
 sg13g2_nand3b_1 _2643_ (.B(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .C(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .Y(_0914_),
    .A_N(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ));
 sg13g2_and2_1 _2644_ (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .B(_0914_),
    .X(_0915_));
 sg13g2_nand3b_1 _2645_ (.B(_0440_),
    .C(_0913_),
    .Y(_0916_),
    .A_N(_0915_));
 sg13g2_nor2_2 _2646_ (.A(net913),
    .B(net973),
    .Y(_0917_));
 sg13g2_o21ai_1 _2647_ (.B1(_0914_),
    .Y(_0918_),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .A2(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ));
 sg13g2_nand2_1 _2648_ (.Y(_0919_),
    .A(_0441_),
    .B(_0917_));
 sg13g2_nor3_1 _2649_ (.A(_0440_),
    .B(_0914_),
    .C(_0917_),
    .Y(_0920_));
 sg13g2_a21oi_1 _2650_ (.A1(_2012_),
    .A2(_0920_),
    .Y(_0921_),
    .B1(_0442_));
 sg13g2_nand3_1 _2651_ (.B(_0919_),
    .C(_0921_),
    .A(_0916_),
    .Y(_0922_));
 sg13g2_nand3_1 _2652_ (.B(net635),
    .C(_0922_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .Y(_0923_));
 sg13g2_nand3_1 _2653_ (.B(net635),
    .C(_0453_),
    .A(net257),
    .Y(_0924_));
 sg13g2_nand2_1 _2654_ (.Y(_0925_),
    .A(net892),
    .B(net703));
 sg13g2_nand3_1 _2655_ (.B(_0924_),
    .C(_0925_),
    .A(_0923_),
    .Y(_0029_));
 sg13g2_nand3_1 _2656_ (.B(_0693_),
    .C(_0743_),
    .A(_0675_),
    .Y(_0926_));
 sg13g2_o21ai_1 _2657_ (.B1(_0926_),
    .Y(_0927_),
    .A1(_0700_),
    .A2(_0769_));
 sg13g2_o21ai_1 _2658_ (.B1(net868),
    .Y(_0928_),
    .A1(_0840_),
    .A2(_0927_));
 sg13g2_nand3_1 _2659_ (.B(net618),
    .C(_0726_),
    .A(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .Y(_0929_));
 sg13g2_o21ai_1 _2660_ (.B1(_0928_),
    .Y(_0002_),
    .A1(_0741_),
    .A2(_0929_));
 sg13g2_o21ai_1 _2661_ (.B1(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .Y(_0930_),
    .A1(_0444_),
    .A2(_0918_));
 sg13g2_o21ai_1 _2662_ (.B1(_0441_),
    .Y(_0931_),
    .A1(_2008_),
    .A2(_2009_));
 sg13g2_nor2_1 _2663_ (.A(_0930_),
    .B(_0931_),
    .Y(_0932_));
 sg13g2_a21o_2 _2664_ (.A2(_0932_),
    .A1(net935),
    .B1(net703),
    .X(_0933_));
 sg13g2_nand2_1 _2665_ (.Y(_0934_),
    .A(_2012_),
    .B(_0450_));
 sg13g2_nand2_1 _2666_ (.Y(_0935_),
    .A(net515),
    .B(_0447_));
 sg13g2_nor2b_1 _2667_ (.A(_0442_),
    .B_N(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .Y(_0936_));
 sg13g2_nand3_1 _2668_ (.B(_0914_),
    .C(_0936_),
    .A(_0441_),
    .Y(_0937_));
 sg13g2_nor2_1 _2669_ (.A(_0917_),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_nand4_1 _2670_ (.B(_0915_),
    .C(_0919_),
    .A(net935),
    .Y(_0939_),
    .D(_0936_));
 sg13g2_inv_1 _2671_ (.Y(_0940_),
    .A(_0939_));
 sg13g2_a221oi_1 _2672_ (.B2(net635),
    .C1(_0940_),
    .B1(_0938_),
    .A1(net1012),
    .Y(_0941_),
    .A2(net579));
 sg13g2_o21ai_1 _2673_ (.B1(_0941_),
    .Y(_0030_),
    .A1(_0934_),
    .A2(_0935_));
 sg13g2_nand2_1 _2674_ (.Y(_0942_),
    .A(net515),
    .B(_0443_));
 sg13g2_o21ai_1 _2675_ (.B1(_0942_),
    .Y(_0943_),
    .A1(net351),
    .A2(_0455_));
 sg13g2_a22oi_1 _2676_ (.Y(_0944_),
    .B1(net635),
    .B2(_0943_),
    .A2(net704),
    .A1(net515));
 sg13g2_inv_1 _2677_ (.Y(_0031_),
    .A(_0944_));
 sg13g2_nand2_1 _2678_ (.Y(_0945_),
    .A(net257),
    .B(net703));
 sg13g2_nand3_1 _2679_ (.B(_0440_),
    .C(net635),
    .A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .Y(_0946_));
 sg13g2_o21ai_1 _2680_ (.B1(_0945_),
    .Y(_0032_),
    .A1(_0913_),
    .A2(_0946_));
 sg13g2_nor2_1 _2681_ (.A(net711),
    .B(_1959_),
    .Y(_0947_));
 sg13g2_nand2_1 _2682_ (.Y(_0948_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .B(_0947_));
 sg13g2_nand3_1 _2683_ (.B(net393),
    .C(net402),
    .A(net740),
    .Y(_0949_));
 sg13g2_nand2_1 _2684_ (.Y(_0950_),
    .A(net342),
    .B(_0949_));
 sg13g2_o21ai_1 _2685_ (.B1(net343),
    .Y(_0033_),
    .A1(_1960_),
    .A2(_0948_));
 sg13g2_a22oi_1 _2686_ (.Y(_0951_),
    .B1(_0948_),
    .B2(net497),
    .A2(_1983_),
    .A1(net740));
 sg13g2_inv_1 _2687_ (.Y(_0034_),
    .A(net498));
 sg13g2_nor2_2 _2688_ (.A(net342),
    .B(net987),
    .Y(_0952_));
 sg13g2_a21oi_1 _2689_ (.A1(_1961_),
    .A2(_0949_),
    .Y(_0035_),
    .B1(_0952_));
 sg13g2_nor2_1 _2690_ (.A(net621),
    .B(_2005_),
    .Y(_0953_));
 sg13g2_nor2_1 _2691_ (.A(net931),
    .B(net556),
    .Y(_0954_));
 sg13g2_a21oi_1 _2692_ (.A1(net623),
    .A2(net705),
    .Y(_0955_),
    .B1(net556));
 sg13g2_nor3_1 _2693_ (.A(_0953_),
    .B(net702),
    .C(net557),
    .Y(_0036_));
 sg13g2_o21ai_1 _2694_ (.B1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .Y(_0956_),
    .A1(net622),
    .A2(_2003_));
 sg13g2_o21ai_1 _2695_ (.B1(_0956_),
    .Y(_0037_),
    .A1(net382),
    .A2(_2000_));
 sg13g2_nand2_1 _2696_ (.Y(_0957_),
    .A(net556),
    .B(_0953_));
 sg13g2_o21ai_1 _2697_ (.B1(net829),
    .Y(_0958_),
    .A1(net622),
    .A2(_2003_));
 sg13g2_nand2_1 _2698_ (.Y(_0038_),
    .A(_0957_),
    .B(net562));
 sg13g2_nand2_1 _2699_ (.Y(_0959_),
    .A(net970),
    .B(_0832_));
 sg13g2_nand3_1 _2700_ (.B(_0713_),
    .C(_0780_),
    .A(_0695_),
    .Y(_0960_));
 sg13g2_nand2_1 _2701_ (.Y(_0003_),
    .A(_0959_),
    .B(_0960_));
 sg13g2_and2_1 _2702_ (.A(net51),
    .B(net48),
    .X(_0041_));
 sg13g2_xnor2_1 _2703_ (.Y(_0961_),
    .A(net810),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ));
 sg13g2_xnor2_1 _2704_ (.Y(_0962_),
    .A(net814),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ));
 sg13g2_xor2_1 _2705_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .A(net806),
    .X(_0963_));
 sg13g2_xnor2_1 _2706_ (.Y(_0964_),
    .A(net807),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ));
 sg13g2_nand3_1 _2707_ (.B(_0962_),
    .C(_0964_),
    .A(_0961_),
    .Y(_0965_));
 sg13g2_o21ai_1 _2708_ (.B1(net735),
    .Y(_0966_),
    .A1(_0963_),
    .A2(_0965_));
 sg13g2_nand2b_1 _2709_ (.Y(_0967_),
    .B(net533),
    .A_N(net11));
 sg13g2_nand2_1 _2710_ (.Y(_0042_),
    .A(_0966_),
    .B(_0967_));
 sg13g2_xnor2_1 _2711_ (.Y(_0968_),
    .A(net386),
    .B(net46));
 sg13g2_xnor2_1 _2712_ (.Y(_0969_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .B(net47));
 sg13g2_nand2_1 _2713_ (.Y(_0970_),
    .A(_0968_),
    .B(_0969_));
 sg13g2_nor2_1 _2714_ (.A(net49),
    .B(_0970_),
    .Y(_0046_));
 sg13g2_nand2b_1 _2715_ (.Y(_0971_),
    .B(net521),
    .A_N(net49));
 sg13g2_a21oi_1 _2716_ (.A1(net704),
    .A2(_0971_),
    .Y(_0047_),
    .B1(_0970_));
 sg13g2_nor2_2 _2717_ (.A(net703),
    .B(_0939_),
    .Y(_0972_));
 sg13g2_nor2_1 _2718_ (.A(net529),
    .B(net599),
    .Y(_0973_));
 sg13g2_nor2_1 _2719_ (.A(net743),
    .B(_0973_),
    .Y(_0045_));
 sg13g2_a21oi_1 _2720_ (.A1(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ),
    .A2(net635),
    .Y(_0974_),
    .B1(net263));
 sg13g2_nor2_1 _2721_ (.A(net741),
    .B(net264),
    .Y(_0044_));
 sg13g2_nor2_1 _2722_ (.A(net519),
    .B(_0454_),
    .Y(_0975_));
 sg13g2_nor2_1 _2723_ (.A(net741),
    .B(net520),
    .Y(_0043_));
 sg13g2_a21oi_2 _2724_ (.B1(_1893_),
    .Y(net38),
    .A2(_1975_),
    .A1(net829));
 sg13g2_a21oi_2 _2725_ (.B1(_0054_),
    .Y(net40),
    .A2(_1975_),
    .A1(net829));
 sg13g2_xor2_1 _2726_ (.B(net48),
    .A(net51),
    .X(_0040_));
 sg13g2_nor2b_1 _2727_ (.A(\u_usb_cdc.bus_reset ),
    .B_N(net722),
    .Y(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ));
 sg13g2_nand2b_1 _2728_ (.Y(_0976_),
    .B(_0601_),
    .A_N(_0469_));
 sg13g2_a21oi_1 _2729_ (.A1(_1902_),
    .A2(_0468_),
    .Y(_0977_),
    .B1(_0466_));
 sg13g2_nand2_1 _2730_ (.Y(_0978_),
    .A(\u_usb_cdc.u_sie.phy_state_q[9] ),
    .B(_0496_));
 sg13g2_o21ai_1 _2731_ (.B1(_0976_),
    .Y(_0979_),
    .A1(_0977_),
    .A2(_0978_));
 sg13g2_a22oi_1 _2732_ (.Y(_0980_),
    .B1(_0979_),
    .B2(_0494_),
    .A2(_0601_),
    .A1(_0498_));
 sg13g2_nor2_1 _2733_ (.A(\u_usb_cdc.u_sie.phy_state_q[8] ),
    .B(net832),
    .Y(_0981_));
 sg13g2_nor4_1 _2734_ (.A(net745),
    .B(_0595_),
    .C(_0599_),
    .D(_0981_),
    .Y(_0982_));
 sg13g2_and2_1 _2735_ (.A(_0980_),
    .B(_0982_),
    .X(_0983_));
 sg13g2_inv_1 _2736_ (.Y(_0984_),
    .A(_0983_));
 sg13g2_nor2b_1 _2737_ (.A(net767),
    .B_N(net169),
    .Y(_0985_));
 sg13g2_a21oi_1 _2738_ (.A1(\u_usb_cdc.endp[0] ),
    .A2(\u_usb_cdc.u_sie.out_toggle_q[1] ),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_xnor2_1 _2739_ (.Y(_0987_),
    .A(\u_usb_cdc.u_sie.pid_q[3] ),
    .B(_0986_));
 sg13g2_nor4_1 _2740_ (.A(\u_usb_cdc.endp[3] ),
    .B(_1985_),
    .C(_0984_),
    .D(_0987_),
    .Y(_0988_));
 sg13g2_a21oi_1 _2741_ (.A1(_1906_),
    .A2(_0988_),
    .Y(_0989_),
    .B1(net169));
 sg13g2_a221oi_1 _2742_ (.B2(_0988_),
    .C1(net170),
    .B1(_0985_),
    .A1(_1903_),
    .Y(_0067_),
    .A2(_0983_));
 sg13g2_nor4_1 _2743_ (.A(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .B(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .C(_0557_),
    .D(_0748_),
    .Y(_0990_));
 sg13g2_nor2_1 _2744_ (.A(net341),
    .B(net271),
    .Y(_0991_));
 sg13g2_nand2_1 _2745_ (.Y(_0992_),
    .A(net518),
    .B(_0991_));
 sg13g2_nor2_1 _2746_ (.A(net423),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_a21oi_1 _2747_ (.A1(_1955_),
    .A2(_0993_),
    .Y(_0994_),
    .B1(net842));
 sg13g2_nor2b_1 _2748_ (.A(_0994_),
    .B_N(_0990_),
    .Y(_0995_));
 sg13g2_nor2_1 _2749_ (.A(net747),
    .B(_0995_),
    .Y(_0996_));
 sg13g2_nand3_1 _2750_ (.B(_0604_),
    .C(_0996_),
    .A(_0590_),
    .Y(_0997_));
 sg13g2_a21oi_1 _2751_ (.A1(net833),
    .A2(_0528_),
    .Y(_0998_),
    .B1(_0997_));
 sg13g2_nand2_1 _2752_ (.Y(_0999_),
    .A(_0594_),
    .B(_0604_));
 sg13g2_nand2b_1 _2753_ (.Y(_1000_),
    .B(net633),
    .A_N(net769));
 sg13g2_nor4_1 _2754_ (.A(_0987_),
    .B(_0998_),
    .C(_0999_),
    .D(_1000_),
    .Y(_1001_));
 sg13g2_xnor2_1 _2755_ (.Y(_1002_),
    .A(net849),
    .B(_1001_));
 sg13g2_a21oi_1 _2756_ (.A1(net739),
    .A2(_0995_),
    .Y(_0068_),
    .B1(net850));
 sg13g2_nand2_1 _2757_ (.Y(_1003_),
    .A(net765),
    .B(_0889_));
 sg13g2_nor2_1 _2758_ (.A(net766),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_o21ai_1 _2759_ (.B1(net745),
    .Y(_1005_),
    .A1(net832),
    .A2(_1004_));
 sg13g2_o21ai_1 _2760_ (.B1(_1005_),
    .Y(_1006_),
    .A1(net836),
    .A2(_0601_));
 sg13g2_nor4_1 _2761_ (.A(net762),
    .B(net1011),
    .C(_1989_),
    .D(_0882_),
    .Y(_1007_));
 sg13g2_nand2_1 _2762_ (.Y(_1008_),
    .A(_1004_),
    .B(_1007_));
 sg13g2_a21oi_1 _2763_ (.A1(net836),
    .A2(_1008_),
    .Y(_1009_),
    .B1(_1006_));
 sg13g2_nand3_1 _2764_ (.B(_0980_),
    .C(_1009_),
    .A(net591),
    .Y(_1010_));
 sg13g2_xnor2_1 _2765_ (.Y(_1011_),
    .A(_1966_),
    .B(net634));
 sg13g2_nor3_1 _2766_ (.A(net832),
    .B(_1010_),
    .C(_1011_),
    .Y(_1012_));
 sg13g2_a21oi_1 _2767_ (.A1(_1966_),
    .A2(_1010_),
    .Y(_0069_),
    .B1(_1012_));
 sg13g2_nand4_1 _2768_ (.B(_0598_),
    .C(_1004_),
    .A(net836),
    .Y(_1013_),
    .D(_1007_));
 sg13g2_and4_1 _2769_ (.A(net836),
    .B(_0598_),
    .C(_1004_),
    .D(_1007_),
    .X(_1014_));
 sg13g2_nand2_1 _2770_ (.Y(_1015_),
    .A(net633),
    .B(_1014_));
 sg13g2_nor4_1 _2771_ (.A(\u_usb_cdc.endp[0] ),
    .B(_1907_),
    .C(\u_usb_cdc.endp[3] ),
    .D(\u_usb_cdc.endp[2] ),
    .Y(_1016_));
 sg13g2_a22oi_1 _2772_ (.Y(_1017_),
    .B1(_1016_),
    .B2(\u_usb_cdc.u_sie.in_toggle_q[2] ),
    .A2(net633),
    .A1(\u_usb_cdc.u_sie.in_toggle_q[1] ));
 sg13g2_o21ai_1 _2773_ (.B1(_1017_),
    .Y(_1018_),
    .A1(_1966_),
    .A2(_0573_));
 sg13g2_a21oi_1 _2774_ (.A1(_1907_),
    .A2(_1987_),
    .Y(_1019_),
    .B1(_1908_));
 sg13g2_nor3_1 _2775_ (.A(_1013_),
    .B(_1018_),
    .C(_1019_),
    .Y(_1020_));
 sg13g2_a22oi_1 _2776_ (.Y(_1021_),
    .B1(_1020_),
    .B2(_0574_),
    .A2(_1015_),
    .A1(net923));
 sg13g2_a21o_1 _2777_ (.A2(_0993_),
    .A1(net479),
    .B1(net842),
    .X(_1022_));
 sg13g2_and2_1 _2778_ (.A(net739),
    .B(_0990_),
    .X(_1023_));
 sg13g2_a21oi_1 _2779_ (.A1(_1022_),
    .A2(_1023_),
    .Y(_0070_),
    .B1(net924));
 sg13g2_nand2_1 _2780_ (.Y(_1024_),
    .A(_1014_),
    .B(_1016_));
 sg13g2_nand2_1 _2781_ (.Y(_1025_),
    .A(net354),
    .B(_1024_));
 sg13g2_nand3_1 _2782_ (.B(_1987_),
    .C(_1020_),
    .A(\u_usb_cdc.endp[1] ),
    .Y(_1026_));
 sg13g2_nand3_1 _2783_ (.B(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .C(_0991_),
    .A(\u_usb_cdc.u_ctrl_endp.endp_q[1] ),
    .Y(_1027_));
 sg13g2_o21ai_1 _2784_ (.B1(_1932_),
    .Y(_1028_),
    .A1(\u_usb_cdc.u_ctrl_endp.endp_q[0] ),
    .A2(_1027_));
 sg13g2_a22oi_1 _2785_ (.Y(_0071_),
    .B1(_1028_),
    .B2(_1023_),
    .A2(_1026_),
    .A1(net355));
 sg13g2_nor2_1 _2786_ (.A(\u_usb_cdc.addr[0] ),
    .B(_0870_),
    .Y(_1029_));
 sg13g2_nand2_1 _2787_ (.Y(_1030_),
    .A(net218),
    .B(_0600_));
 sg13g2_a21oi_1 _2788_ (.A1(net761),
    .A2(_0870_),
    .Y(_1031_),
    .B1(_1029_));
 sg13g2_o21ai_1 _2789_ (.B1(net219),
    .Y(_0072_),
    .A1(_0600_),
    .A2(_1031_));
 sg13g2_nand2_1 _2790_ (.Y(_1032_),
    .A(net308),
    .B(net713));
 sg13g2_nor2_1 _2791_ (.A(net829),
    .B(_1993_),
    .Y(_1033_));
 sg13g2_nand2b_2 _2792_ (.Y(_1034_),
    .B(net702),
    .A_N(net829));
 sg13g2_a221oi_1 _2793_ (.B2(net702),
    .C1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .B1(_1994_),
    .A1(_1893_),
    .Y(_1035_),
    .A2(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ));
 sg13g2_a21oi_1 _2794_ (.A1(_2006_),
    .A2(_1035_),
    .Y(_1036_),
    .B1(_1996_));
 sg13g2_a22oi_1 _2795_ (.Y(_1037_),
    .B1(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .B2(net623),
    .A2(net743),
    .A1(_1893_));
 sg13g2_o21ai_1 _2796_ (.B1(_1032_),
    .Y(_0073_),
    .A1(_1036_),
    .A2(_1037_));
 sg13g2_nand2_1 _2797_ (.Y(_1038_),
    .A(net941),
    .B(net10));
 sg13g2_nor2_1 _2798_ (.A(net827),
    .B(net825),
    .Y(_1039_));
 sg13g2_nor3_2 _2799_ (.A(net828),
    .B(net827),
    .C(net824),
    .Y(_1040_));
 sg13g2_a21oi_1 _2800_ (.A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .A2(_1039_),
    .Y(_1041_),
    .B1(net997));
 sg13g2_xnor2_1 _2801_ (.Y(_1042_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .B(_1041_));
 sg13g2_nand2_2 _2802_ (.Y(_1043_),
    .A(net828),
    .B(net827));
 sg13g2_nand4_1 _2803_ (.B(net1066),
    .C(net824),
    .A(net828),
    .Y(_1044_),
    .D(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ));
 sg13g2_xor2_1 _2804_ (.B(net1053),
    .A(net997),
    .X(_1045_));
 sg13g2_xnor2_1 _2805_ (.Y(_1046_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .B(_1045_));
 sg13g2_nand2b_1 _2806_ (.Y(_1047_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .A_N(_1040_));
 sg13g2_o21ai_1 _2807_ (.B1(_1047_),
    .Y(_1048_),
    .A1(net707),
    .A2(_1043_));
 sg13g2_xnor2_1 _2808_ (.Y(_1049_),
    .A(net825),
    .B(_1043_));
 sg13g2_xnor2_1 _2809_ (.Y(_1050_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .B(_1049_));
 sg13g2_nand4_1 _2810_ (.B(_1044_),
    .C(_1046_),
    .A(_1042_),
    .Y(_1051_),
    .D(_1050_));
 sg13g2_and2_1 _2811_ (.A(_1044_),
    .B(_1048_),
    .X(_1052_));
 sg13g2_xor2_1 _2812_ (.B(_1052_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .X(_1053_));
 sg13g2_o21ai_1 _2813_ (.B1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ),
    .Y(_1054_),
    .A1(_1051_),
    .A2(_1053_));
 sg13g2_or2_1 _2814_ (.X(_1055_),
    .B(_1054_),
    .A(net714));
 sg13g2_nand2_2 _2815_ (.Y(_1056_),
    .A(net542),
    .B(_1055_));
 sg13g2_nand2_1 _2816_ (.Y(_0074_),
    .A(net638),
    .B(_1056_));
 sg13g2_mux2_1 _2817_ (.A0(net2),
    .A1(net1022),
    .S(net637),
    .X(_0075_));
 sg13g2_mux2_1 _2818_ (.A0(net3),
    .A1(net1021),
    .S(net637),
    .X(_0076_));
 sg13g2_mux2_1 _2819_ (.A0(net4),
    .A1(net1032),
    .S(net637),
    .X(_0077_));
 sg13g2_mux2_1 _2820_ (.A0(net5),
    .A1(net1040),
    .S(net637),
    .X(_0078_));
 sg13g2_mux2_1 _2821_ (.A0(net6),
    .A1(net1033),
    .S(net637),
    .X(_0079_));
 sg13g2_mux2_1 _2822_ (.A0(net7),
    .A1(net1041),
    .S(net637),
    .X(_0080_));
 sg13g2_mux2_1 _2823_ (.A0(net8),
    .A1(net1042),
    .S(net637),
    .X(_0081_));
 sg13g2_mux2_1 _2824_ (.A0(net9),
    .A1(net1039),
    .S(net637),
    .X(_0082_));
 sg13g2_nor2_2 _2825_ (.A(net714),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .Y(_1057_));
 sg13g2_nand2_2 _2826_ (.Y(_1058_),
    .A(_1040_),
    .B(_1057_));
 sg13g2_mux2_1 _2827_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .A1(net378),
    .S(_1058_),
    .X(_0083_));
 sg13g2_mux2_1 _2828_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .A1(net442),
    .S(_1058_),
    .X(_0084_));
 sg13g2_mux2_1 _2829_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .A1(net424),
    .S(_1058_),
    .X(_0085_));
 sg13g2_mux2_1 _2830_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .A1(net407),
    .S(_1058_),
    .X(_0086_));
 sg13g2_mux2_1 _2831_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .A1(net397),
    .S(_1058_),
    .X(_0087_));
 sg13g2_mux2_1 _2832_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .A1(net554),
    .S(_1058_),
    .X(_0088_));
 sg13g2_mux2_1 _2833_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .A1(net380),
    .S(_1058_),
    .X(_0089_));
 sg13g2_mux2_1 _2834_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .A1(net438),
    .S(_1058_),
    .X(_0090_));
 sg13g2_nand3_1 _2835_ (.B(_1039_),
    .C(_1057_),
    .A(net828),
    .Y(_1059_));
 sg13g2_nand2_1 _2836_ (.Y(_1060_),
    .A(net95),
    .B(_1059_));
 sg13g2_nor2b_2 _2837_ (.A(net827),
    .B_N(net828),
    .Y(_1061_));
 sg13g2_nand2_1 _2838_ (.Y(_1062_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .B(net636));
 sg13g2_xnor2_1 _2839_ (.Y(_1063_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .B(_1040_));
 sg13g2_nand3_1 _2840_ (.B(net707),
    .C(_1063_),
    .A(net736),
    .Y(_1064_));
 sg13g2_o21ai_1 _2841_ (.B1(_1060_),
    .Y(_0091_),
    .A1(_1062_),
    .A2(net616));
 sg13g2_nand2_1 _2842_ (.Y(_1065_),
    .A(net75),
    .B(_1059_));
 sg13g2_nand2_1 _2843_ (.Y(_1066_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .B(net636));
 sg13g2_o21ai_1 _2844_ (.B1(_1065_),
    .Y(_0092_),
    .A1(net616),
    .A2(_1066_));
 sg13g2_nand2_1 _2845_ (.Y(_1067_),
    .A(net191),
    .B(_1059_));
 sg13g2_nand2_1 _2846_ (.Y(_1068_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .B(net636));
 sg13g2_o21ai_1 _2847_ (.B1(_1067_),
    .Y(_0093_),
    .A1(net616),
    .A2(_1068_));
 sg13g2_nand2_1 _2848_ (.Y(_1069_),
    .A(net137),
    .B(_1059_));
 sg13g2_nand2_1 _2849_ (.Y(_1070_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .B(net636));
 sg13g2_o21ai_1 _2850_ (.B1(_1069_),
    .Y(_0094_),
    .A1(net616),
    .A2(_1070_));
 sg13g2_nand2_1 _2851_ (.Y(_1071_),
    .A(net69),
    .B(_1059_));
 sg13g2_nand2_1 _2852_ (.Y(_1072_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .B(net636));
 sg13g2_o21ai_1 _2853_ (.B1(_1071_),
    .Y(_0095_),
    .A1(net616),
    .A2(_1072_));
 sg13g2_nand2_1 _2854_ (.Y(_1073_),
    .A(net253),
    .B(_1059_));
 sg13g2_nand2_1 _2855_ (.Y(_1074_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .B(net636));
 sg13g2_o21ai_1 _2856_ (.B1(_1073_),
    .Y(_0096_),
    .A1(net616),
    .A2(_1074_));
 sg13g2_nand2_1 _2857_ (.Y(_1075_),
    .A(net151),
    .B(_1059_));
 sg13g2_nand2_1 _2858_ (.Y(_1076_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .B(net636));
 sg13g2_o21ai_1 _2859_ (.B1(_1075_),
    .Y(_0097_),
    .A1(_1064_),
    .A2(_1076_));
 sg13g2_nand2_1 _2860_ (.Y(_1077_),
    .A(net91),
    .B(_1059_));
 sg13g2_nand2_1 _2861_ (.Y(_1078_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .B(net636));
 sg13g2_o21ai_1 _2862_ (.B1(_1077_),
    .Y(_0098_),
    .A1(_1064_),
    .A2(_1078_));
 sg13g2_nor2b_2 _2863_ (.A(net828),
    .B_N(net827),
    .Y(_1079_));
 sg13g2_nand2b_2 _2864_ (.Y(_1080_),
    .B(_1079_),
    .A_N(net616));
 sg13g2_nand2_1 _2865_ (.Y(_1081_),
    .A(net162),
    .B(_1080_));
 sg13g2_and3_2 _2866_ (.X(_1082_),
    .A(net736),
    .B(_1063_),
    .C(_1079_));
 sg13g2_nand2_1 _2867_ (.Y(_1083_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2868_ (.B1(_1081_),
    .Y(_0099_),
    .A1(net826),
    .A2(_1083_));
 sg13g2_nand2_1 _2869_ (.Y(_1084_),
    .A(net89),
    .B(_1080_));
 sg13g2_nand2_1 _2870_ (.Y(_1085_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2871_ (.B1(_1084_),
    .Y(_0100_),
    .A1(net826),
    .A2(_1085_));
 sg13g2_nand2_1 _2872_ (.Y(_1086_),
    .A(net178),
    .B(_1080_));
 sg13g2_nand2_1 _2873_ (.Y(_1087_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2874_ (.B1(_1086_),
    .Y(_0101_),
    .A1(net826),
    .A2(_1087_));
 sg13g2_nand2_1 _2875_ (.Y(_1088_),
    .A(net184),
    .B(_1080_));
 sg13g2_nand2_1 _2876_ (.Y(_1089_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2877_ (.B1(_1088_),
    .Y(_0102_),
    .A1(net826),
    .A2(_1089_));
 sg13g2_nand2_1 _2878_ (.Y(_1090_),
    .A(net61),
    .B(_1080_));
 sg13g2_nand2_1 _2879_ (.Y(_1091_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2880_ (.B1(_1090_),
    .Y(_0103_),
    .A1(net824),
    .A2(_1091_));
 sg13g2_nand2_1 _2881_ (.Y(_1092_),
    .A(net93),
    .B(_1080_));
 sg13g2_nand2_1 _2882_ (.Y(_1093_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2883_ (.B1(_1092_),
    .Y(_0104_),
    .A1(net826),
    .A2(_1093_));
 sg13g2_nand2_1 _2884_ (.Y(_1094_),
    .A(net147),
    .B(_1080_));
 sg13g2_nand2_1 _2885_ (.Y(_1095_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2886_ (.B1(_1094_),
    .Y(_0105_),
    .A1(net824),
    .A2(_1095_));
 sg13g2_nand2_1 _2887_ (.Y(_1096_),
    .A(net67),
    .B(_1080_));
 sg13g2_nand2_1 _2888_ (.Y(_1097_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .B(_1082_));
 sg13g2_o21ai_1 _2889_ (.B1(_1096_),
    .Y(_0106_),
    .A1(net824),
    .A2(_1097_));
 sg13g2_or2_1 _2890_ (.X(_1098_),
    .B(net616),
    .A(_1043_));
 sg13g2_mux2_1 _2891_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .A1(net418),
    .S(_1098_),
    .X(_0107_));
 sg13g2_mux2_1 _2892_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .A1(net489),
    .S(_1098_),
    .X(_0108_));
 sg13g2_mux2_1 _2893_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .A1(net426),
    .S(_1098_),
    .X(_0109_));
 sg13g2_mux2_1 _2894_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .A1(net452),
    .S(_1098_),
    .X(_0110_));
 sg13g2_mux2_1 _2895_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .A1(net481),
    .S(_1098_),
    .X(_0111_));
 sg13g2_mux2_1 _2896_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .A1(net410),
    .S(_1098_),
    .X(_0112_));
 sg13g2_mux2_1 _2897_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .A1(net456),
    .S(_1098_),
    .X(_0113_));
 sg13g2_mux2_1 _2898_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .A1(net473),
    .S(_1098_),
    .X(_0114_));
 sg13g2_nand2_2 _2899_ (.Y(_1099_),
    .A(net824),
    .B(_1057_));
 sg13g2_nor3_2 _2900_ (.A(net828),
    .B(net827),
    .C(net615),
    .Y(_1100_));
 sg13g2_mux2_1 _2901_ (.A0(net436),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .S(_1100_),
    .X(_0115_));
 sg13g2_mux2_1 _2902_ (.A0(net471),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .S(_1100_),
    .X(_0116_));
 sg13g2_mux2_1 _2903_ (.A0(net446),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .S(_1100_),
    .X(_0117_));
 sg13g2_mux2_1 _2904_ (.A0(net454),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .S(_1100_),
    .X(_0118_));
 sg13g2_mux2_1 _2905_ (.A0(net467),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .S(_1100_),
    .X(_0119_));
 sg13g2_mux2_1 _2906_ (.A0(net513),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .S(_1100_),
    .X(_0120_));
 sg13g2_mux2_1 _2907_ (.A0(net475),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .S(_1100_),
    .X(_0121_));
 sg13g2_mux2_1 _2908_ (.A0(net376),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .S(_1100_),
    .X(_0122_));
 sg13g2_nand3_1 _2909_ (.B(_1057_),
    .C(_1061_),
    .A(net824),
    .Y(_1101_));
 sg13g2_nand2_1 _2910_ (.Y(_1102_),
    .A(net83),
    .B(_1101_));
 sg13g2_o21ai_1 _2911_ (.B1(_1102_),
    .Y(_0123_),
    .A1(_1062_),
    .A2(net615));
 sg13g2_nand2_1 _2912_ (.Y(_1103_),
    .A(net73),
    .B(_1101_));
 sg13g2_o21ai_1 _2913_ (.B1(_1103_),
    .Y(_0124_),
    .A1(_1066_),
    .A2(net615));
 sg13g2_nand2_1 _2914_ (.Y(_1104_),
    .A(net110),
    .B(_1101_));
 sg13g2_o21ai_1 _2915_ (.B1(_1104_),
    .Y(_0125_),
    .A1(_1068_),
    .A2(net615));
 sg13g2_nand2_1 _2916_ (.Y(_1105_),
    .A(net149),
    .B(_1101_));
 sg13g2_o21ai_1 _2917_ (.B1(_1105_),
    .Y(_0126_),
    .A1(_1070_),
    .A2(net615));
 sg13g2_nand2_1 _2918_ (.Y(_1106_),
    .A(net130),
    .B(_1101_));
 sg13g2_o21ai_1 _2919_ (.B1(_1106_),
    .Y(_0127_),
    .A1(_1072_),
    .A2(net615));
 sg13g2_nand2_1 _2920_ (.Y(_1107_),
    .A(net56),
    .B(_1101_));
 sg13g2_o21ai_1 _2921_ (.B1(_1107_),
    .Y(_0128_),
    .A1(_1074_),
    .A2(net615));
 sg13g2_nand2_1 _2922_ (.Y(_1108_),
    .A(net71),
    .B(_1101_));
 sg13g2_o21ai_1 _2923_ (.B1(_1108_),
    .Y(_0129_),
    .A1(_1076_),
    .A2(_1099_));
 sg13g2_nand2_1 _2924_ (.Y(_1109_),
    .A(net80),
    .B(_1101_));
 sg13g2_o21ai_1 _2925_ (.B1(_1109_),
    .Y(_0130_),
    .A1(_1078_),
    .A2(_1099_));
 sg13g2_nand3_1 _2926_ (.B(_1057_),
    .C(_1079_),
    .A(net824),
    .Y(_1110_));
 sg13g2_nand2_1 _2927_ (.Y(_1111_),
    .A(net155),
    .B(_1110_));
 sg13g2_o21ai_1 _2928_ (.B1(_1111_),
    .Y(_0131_),
    .A1(net707),
    .A2(_1083_));
 sg13g2_nand2_1 _2929_ (.Y(_1112_),
    .A(net114),
    .B(_1110_));
 sg13g2_o21ai_1 _2930_ (.B1(_1112_),
    .Y(_0132_),
    .A1(net707),
    .A2(_1085_));
 sg13g2_nand2_1 _2931_ (.Y(_1113_),
    .A(net124),
    .B(_1110_));
 sg13g2_o21ai_1 _2932_ (.B1(_1113_),
    .Y(_0133_),
    .A1(net707),
    .A2(_1087_));
 sg13g2_nand2_1 _2933_ (.Y(_1114_),
    .A(net159),
    .B(_1110_));
 sg13g2_o21ai_1 _2934_ (.B1(_1114_),
    .Y(_0134_),
    .A1(net707),
    .A2(_1089_));
 sg13g2_nand2_1 _2935_ (.Y(_1115_),
    .A(net126),
    .B(_1110_));
 sg13g2_o21ai_1 _2936_ (.B1(_1115_),
    .Y(_0135_),
    .A1(net707),
    .A2(_1091_));
 sg13g2_nand2_1 _2937_ (.Y(_1116_),
    .A(net106),
    .B(_1110_));
 sg13g2_o21ai_1 _2938_ (.B1(_1116_),
    .Y(_0136_),
    .A1(net707),
    .A2(_1093_));
 sg13g2_nand2_1 _2939_ (.Y(_1117_),
    .A(net87),
    .B(_1110_));
 sg13g2_o21ai_1 _2940_ (.B1(_1117_),
    .Y(_0137_),
    .A1(_1965_),
    .A2(_1095_));
 sg13g2_nand2_1 _2941_ (.Y(_1118_),
    .A(net59),
    .B(_1110_));
 sg13g2_o21ai_1 _2942_ (.B1(_1118_),
    .Y(_0138_),
    .A1(_1965_),
    .A2(_1097_));
 sg13g2_nor2_2 _2943_ (.A(_1043_),
    .B(net615),
    .Y(_1119_));
 sg13g2_mux2_1 _2944_ (.A0(net395),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .S(net603),
    .X(_0139_));
 sg13g2_mux2_1 _2945_ (.A0(net434),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .S(net603),
    .X(_0140_));
 sg13g2_mux2_1 _2946_ (.A0(net511),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .S(net603),
    .X(_0141_));
 sg13g2_mux2_1 _2947_ (.A0(net493),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .S(net603),
    .X(_0142_));
 sg13g2_mux2_1 _2948_ (.A0(net487),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .S(_1119_),
    .X(_0143_));
 sg13g2_mux2_1 _2949_ (.A0(net483),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .S(net603),
    .X(_0144_));
 sg13g2_mux2_1 _2950_ (.A0(net462),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .S(net603),
    .X(_0145_));
 sg13g2_nand2_1 _2951_ (.Y(_1120_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .B(net603));
 sg13g2_o21ai_1 _2952_ (.B1(_1120_),
    .Y(_0146_),
    .A1(_1974_),
    .A2(net603));
 sg13g2_and3_2 _2953_ (.X(_1121_),
    .A(net736),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .C(_1040_));
 sg13g2_mux2_1 _2954_ (.A0(net450),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .S(_1121_),
    .X(_0147_));
 sg13g2_mux2_1 _2955_ (.A0(net430),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .S(_1121_),
    .X(_0148_));
 sg13g2_mux2_1 _2956_ (.A0(net464),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .S(_1121_),
    .X(_0149_));
 sg13g2_mux2_1 _2957_ (.A0(net477),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .S(_1121_),
    .X(_0150_));
 sg13g2_mux2_1 _2958_ (.A0(net448),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .S(_1121_),
    .X(_0151_));
 sg13g2_mux2_1 _2959_ (.A0(net432),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .S(_1121_),
    .X(_0152_));
 sg13g2_mux2_1 _2960_ (.A0(net469),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .S(_1121_),
    .X(_0153_));
 sg13g2_mux2_1 _2961_ (.A0(net491),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .S(_1121_),
    .X(_0154_));
 sg13g2_nand2_1 _2962_ (.Y(_1122_),
    .A(net739),
    .B(net632));
 sg13g2_a21oi_2 _2963_ (.B1(_1122_),
    .Y(_1123_),
    .A2(_0621_),
    .A1(_0620_));
 sg13g2_mux2_1 _2964_ (.A0(_1045_),
    .A1(net827),
    .S(_1054_),
    .X(_1124_));
 sg13g2_mux2_1 _2965_ (.A0(net870),
    .A1(_1124_),
    .S(_1123_),
    .X(_0155_));
 sg13g2_mux2_1 _2966_ (.A0(_1049_),
    .A1(net825),
    .S(_1054_),
    .X(_1125_));
 sg13g2_mux2_1 _2967_ (.A0(net857),
    .A1(_1125_),
    .S(_1123_),
    .X(_0156_));
 sg13g2_mux2_1 _2968_ (.A0(_1052_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .S(_1054_),
    .X(_1126_));
 sg13g2_mux2_1 _2969_ (.A0(net901),
    .A1(_1126_),
    .S(_1123_),
    .X(_0157_));
 sg13g2_o21ai_1 _2970_ (.B1(net638),
    .Y(_1127_),
    .A1(net941),
    .A2(_1056_));
 sg13g2_inv_1 _2971_ (.Y(_0158_),
    .A(_1127_));
 sg13g2_mux2_1 _2972_ (.A0(_1041_),
    .A1(net997),
    .S(_1055_),
    .X(_0159_));
 sg13g2_mux2_1 _2973_ (.A0(_1045_),
    .A1(net827),
    .S(_1055_),
    .X(_0160_));
 sg13g2_mux2_1 _2974_ (.A0(_1049_),
    .A1(net825),
    .S(_1055_),
    .X(_0161_));
 sg13g2_mux2_1 _2975_ (.A0(_1052_),
    .A1(net1020),
    .S(_1055_),
    .X(_0162_));
 sg13g2_nand2_2 _2976_ (.Y(_1128_),
    .A(\u_usb_cdc.sie_in_req ),
    .B(net631));
 sg13g2_nand2_1 _2977_ (.Y(_1129_),
    .A(net1034),
    .B(_1128_));
 sg13g2_nand3_1 _2978_ (.B(_1123_),
    .C(_1128_),
    .A(\u_usb_cdc.sie_in_data_ack ),
    .Y(_1130_));
 sg13g2_nand2_1 _2979_ (.Y(_1131_),
    .A(net301),
    .B(_1130_));
 sg13g2_o21ai_1 _2980_ (.B1(_1131_),
    .Y(_0163_),
    .A1(_1912_),
    .A2(_1130_));
 sg13g2_mux2_1 _2981_ (.A0(net794),
    .A1(net927),
    .S(_1130_),
    .X(_0164_));
 sg13g2_nand2_1 _2982_ (.Y(_1132_),
    .A(net280),
    .B(_1130_));
 sg13g2_o21ai_1 _2983_ (.B1(_1132_),
    .Y(_0165_),
    .A1(_1913_),
    .A2(_1130_));
 sg13g2_nand2_1 _2984_ (.Y(_1133_),
    .A(net335),
    .B(_1130_));
 sg13g2_o21ai_1 _2985_ (.B1(_1133_),
    .Y(_0166_),
    .A1(_1914_),
    .A2(_1130_));
 sg13g2_nor2_2 _2986_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .Y(_1134_));
 sg13g2_nand2_2 _2987_ (.Y(_1135_),
    .A(net709),
    .B(_1134_));
 sg13g2_nor2_2 _2988_ (.A(net714),
    .B(net822),
    .Y(_1136_));
 sg13g2_nand2b_2 _2989_ (.Y(_1137_),
    .B(_1136_),
    .A_N(net630));
 sg13g2_nand2_1 _2990_ (.Y(_1138_),
    .A(net255),
    .B(net613));
 sg13g2_o21ai_1 _2991_ (.B1(_1138_),
    .Y(_0167_),
    .A1(net721),
    .A2(_1137_));
 sg13g2_nand2_1 _2992_ (.Y(_1139_),
    .A(net97),
    .B(net613));
 sg13g2_o21ai_1 _2993_ (.B1(_1139_),
    .Y(_0168_),
    .A1(net720),
    .A2(net613));
 sg13g2_nand2_1 _2994_ (.Y(_1140_),
    .A(net82),
    .B(net614));
 sg13g2_o21ai_1 _2995_ (.B1(_1140_),
    .Y(_0169_),
    .A1(net718),
    .A2(net614));
 sg13g2_nand2_1 _2996_ (.Y(_1141_),
    .A(net63),
    .B(net614));
 sg13g2_o21ai_1 _2997_ (.B1(_1141_),
    .Y(_0170_),
    .A1(net719),
    .A2(net614));
 sg13g2_nand2_1 _2998_ (.Y(_1142_),
    .A(net157),
    .B(net614));
 sg13g2_o21ai_1 _2999_ (.B1(_1142_),
    .Y(_0171_),
    .A1(_1899_),
    .A2(net613));
 sg13g2_nand2_1 _3000_ (.Y(_1143_),
    .A(net232),
    .B(net613));
 sg13g2_o21ai_1 _3001_ (.B1(_1143_),
    .Y(_0172_),
    .A1(_1898_),
    .A2(net613));
 sg13g2_nand2_1 _3002_ (.Y(_1144_),
    .A(net54),
    .B(net614));
 sg13g2_o21ai_1 _3003_ (.B1(_1144_),
    .Y(_0173_),
    .A1(_1901_),
    .A2(net614));
 sg13g2_nand2_1 _3004_ (.Y(_1145_),
    .A(net229),
    .B(net613));
 sg13g2_o21ai_1 _3005_ (.B1(_1145_),
    .Y(_0174_),
    .A1(net717),
    .A2(net613));
 sg13g2_nand4_1 _3006_ (.B(net823),
    .C(net709),
    .A(net735),
    .Y(_1146_),
    .D(_1134_));
 sg13g2_nand2_1 _3007_ (.Y(_1147_),
    .A(net104),
    .B(_1146_));
 sg13g2_nor3_2 _3008_ (.A(net822),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .C(net820),
    .Y(_1148_));
 sg13g2_xnor2_1 _3009_ (.Y(_1149_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .B(_1148_));
 sg13g2_and3_2 _3010_ (.X(_1150_),
    .A(net735),
    .B(_1962_),
    .C(_1149_));
 sg13g2_nand3_1 _3011_ (.B(net823),
    .C(_1150_),
    .A(net761),
    .Y(_1151_));
 sg13g2_o21ai_1 _3012_ (.B1(_1147_),
    .Y(_0175_),
    .A1(net821),
    .A2(_1151_));
 sg13g2_nand2_1 _3013_ (.Y(_1152_),
    .A(net216),
    .B(_1146_));
 sg13g2_nand3_1 _3014_ (.B(net823),
    .C(_1150_),
    .A(net759),
    .Y(_1153_));
 sg13g2_o21ai_1 _3015_ (.B1(_1152_),
    .Y(_0176_),
    .A1(net821),
    .A2(_1153_));
 sg13g2_nand2_1 _3016_ (.Y(_1154_),
    .A(net122),
    .B(_1146_));
 sg13g2_nand3_1 _3017_ (.B(net823),
    .C(_1150_),
    .A(net756),
    .Y(_1155_));
 sg13g2_o21ai_1 _3018_ (.B1(_1154_),
    .Y(_0177_),
    .A1(net821),
    .A2(_1155_));
 sg13g2_nand2_1 _3019_ (.Y(_1156_),
    .A(net102),
    .B(_1146_));
 sg13g2_nand3_1 _3020_ (.B(net823),
    .C(_1150_),
    .A(net755),
    .Y(_1157_));
 sg13g2_o21ai_1 _3021_ (.B1(_1156_),
    .Y(_0178_),
    .A1(net821),
    .A2(_1157_));
 sg13g2_nand2_1 _3022_ (.Y(_1158_),
    .A(net153),
    .B(_1146_));
 sg13g2_nand3_1 _3023_ (.B(net823),
    .C(_1150_),
    .A(net754),
    .Y(_1159_));
 sg13g2_o21ai_1 _3024_ (.B1(_1158_),
    .Y(_0179_),
    .A1(net821),
    .A2(_1159_));
 sg13g2_nand2_1 _3025_ (.Y(_1160_),
    .A(net225),
    .B(_1146_));
 sg13g2_nand3_1 _3026_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .C(_1150_),
    .A(net753),
    .Y(_1161_));
 sg13g2_o21ai_1 _3027_ (.B1(_1160_),
    .Y(_0180_),
    .A1(net821),
    .A2(_1161_));
 sg13g2_nand2_1 _3028_ (.Y(_1162_),
    .A(net180),
    .B(_1146_));
 sg13g2_nand3_1 _3029_ (.B(net823),
    .C(_1150_),
    .A(net752),
    .Y(_1163_));
 sg13g2_o21ai_1 _3030_ (.B1(_1162_),
    .Y(_0181_),
    .A1(net821),
    .A2(_1163_));
 sg13g2_nand2_1 _3031_ (.Y(_1164_),
    .A(net221),
    .B(_1146_));
 sg13g2_nand3_1 _3032_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .C(_1150_),
    .A(net751),
    .Y(_1165_));
 sg13g2_o21ai_1 _3033_ (.B1(_1164_),
    .Y(_0182_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .A2(_1165_));
 sg13g2_and4_1 _3034_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .B(net709),
    .C(_1964_),
    .D(_1136_),
    .X(_1166_));
 sg13g2_nor2_1 _3035_ (.A(net389),
    .B(net611),
    .Y(_1167_));
 sg13g2_nand2_2 _3036_ (.Y(_1168_),
    .A(net761),
    .B(net630));
 sg13g2_a21oi_1 _3037_ (.A1(net611),
    .A2(_1168_),
    .Y(_0183_),
    .B1(_1167_));
 sg13g2_nor2_1 _3038_ (.A(net546),
    .B(net611),
    .Y(_1169_));
 sg13g2_nand2_2 _3039_ (.Y(_1170_),
    .A(net759),
    .B(net630));
 sg13g2_a21oi_1 _3040_ (.A1(net611),
    .A2(_1170_),
    .Y(_0184_),
    .B1(_1169_));
 sg13g2_nor2_1 _3041_ (.A(net321),
    .B(net611),
    .Y(_1171_));
 sg13g2_nand2_2 _3042_ (.Y(_1172_),
    .A(net756),
    .B(net630));
 sg13g2_a21oi_1 _3043_ (.A1(net611),
    .A2(_1172_),
    .Y(_0185_),
    .B1(_1171_));
 sg13g2_nand2_1 _3044_ (.Y(_1173_),
    .A(net755),
    .B(net630));
 sg13g2_nor2_1 _3045_ (.A(net440),
    .B(net611),
    .Y(_1174_));
 sg13g2_a21oi_1 _3046_ (.A1(net611),
    .A2(_1173_),
    .Y(_0186_),
    .B1(_1174_));
 sg13g2_nor2_1 _3047_ (.A(net299),
    .B(net612),
    .Y(_1175_));
 sg13g2_nand2_2 _3048_ (.Y(_1176_),
    .A(net754),
    .B(net630));
 sg13g2_a21oi_1 _3049_ (.A1(net612),
    .A2(_1176_),
    .Y(_0187_),
    .B1(_1175_));
 sg13g2_nor2_1 _3050_ (.A(net283),
    .B(net612),
    .Y(_1177_));
 sg13g2_nand2_2 _3051_ (.Y(_1178_),
    .A(net753),
    .B(net630));
 sg13g2_a21oi_1 _3052_ (.A1(net612),
    .A2(_1178_),
    .Y(_0188_),
    .B1(_1177_));
 sg13g2_nor2_1 _3053_ (.A(net267),
    .B(net612),
    .Y(_1179_));
 sg13g2_nand2_2 _3054_ (.Y(_1180_),
    .A(net752),
    .B(net630));
 sg13g2_a21oi_1 _3055_ (.A1(net612),
    .A2(_1180_),
    .Y(_0189_),
    .B1(_1179_));
 sg13g2_nor2_1 _3056_ (.A(net314),
    .B(net612),
    .Y(_1181_));
 sg13g2_nand2_2 _3057_ (.Y(_1182_),
    .A(net751),
    .B(_1135_));
 sg13g2_a21oi_1 _3058_ (.A1(net612),
    .A2(_1182_),
    .Y(_0190_),
    .B1(_1181_));
 sg13g2_and2_1 _3059_ (.A(net822),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .X(_1183_));
 sg13g2_nand4_1 _3060_ (.B(net708),
    .C(_1149_),
    .A(net735),
    .Y(_1184_),
    .D(_1183_));
 sg13g2_nand2_1 _3061_ (.Y(_1185_),
    .A(net227),
    .B(net608));
 sg13g2_o21ai_1 _3062_ (.B1(_1185_),
    .Y(_0191_),
    .A1(net721),
    .A2(net608));
 sg13g2_nand2_1 _3063_ (.Y(_1186_),
    .A(net239),
    .B(net608));
 sg13g2_o21ai_1 _3064_ (.B1(_1186_),
    .Y(_0192_),
    .A1(net720),
    .A2(net608));
 sg13g2_nand2_1 _3065_ (.Y(_1187_),
    .A(net66),
    .B(net608));
 sg13g2_o21ai_1 _3066_ (.B1(_1187_),
    .Y(_0193_),
    .A1(net718),
    .A2(net608));
 sg13g2_nand2_1 _3067_ (.Y(_1188_),
    .A(net58),
    .B(net610));
 sg13g2_o21ai_1 _3068_ (.B1(_1188_),
    .Y(_0194_),
    .A1(net719),
    .A2(net610));
 sg13g2_nand2_1 _3069_ (.Y(_1189_),
    .A(net176),
    .B(net609));
 sg13g2_o21ai_1 _3070_ (.B1(_1189_),
    .Y(_0195_),
    .A1(_1899_),
    .A2(net609));
 sg13g2_nand2_1 _3071_ (.Y(_1190_),
    .A(net204),
    .B(net608));
 sg13g2_o21ai_1 _3072_ (.B1(_1190_),
    .Y(_0196_),
    .A1(_1898_),
    .A2(net608));
 sg13g2_nand2_1 _3073_ (.Y(_1191_),
    .A(net182),
    .B(net610));
 sg13g2_o21ai_1 _3074_ (.B1(_1191_),
    .Y(_0197_),
    .A1(_1901_),
    .A2(net610));
 sg13g2_nand2_1 _3075_ (.Y(_1192_),
    .A(net201),
    .B(net609));
 sg13g2_o21ai_1 _3076_ (.B1(_1192_),
    .Y(_0198_),
    .A1(net717),
    .A2(net609));
 sg13g2_nand3_1 _3077_ (.B(_1134_),
    .C(_1136_),
    .A(net820),
    .Y(_1193_));
 sg13g2_nand2_1 _3078_ (.Y(_1194_),
    .A(net242),
    .B(net606));
 sg13g2_o21ai_1 _3079_ (.B1(_1194_),
    .Y(_0199_),
    .A1(net721),
    .A2(net606));
 sg13g2_nand2_1 _3080_ (.Y(_1195_),
    .A(net188),
    .B(net606));
 sg13g2_o21ai_1 _3081_ (.B1(_1195_),
    .Y(_0200_),
    .A1(net720),
    .A2(net606));
 sg13g2_nand2_1 _3082_ (.Y(_1196_),
    .A(net174),
    .B(net606));
 sg13g2_o21ai_1 _3083_ (.B1(_1196_),
    .Y(_0201_),
    .A1(net718),
    .A2(net606));
 sg13g2_nand2_1 _3084_ (.Y(_1197_),
    .A(net77),
    .B(net607));
 sg13g2_o21ai_1 _3085_ (.B1(_1197_),
    .Y(_0202_),
    .A1(net719),
    .A2(net607));
 sg13g2_nand2_1 _3086_ (.Y(_1198_),
    .A(net240),
    .B(net606));
 sg13g2_o21ai_1 _3087_ (.B1(_1198_),
    .Y(_0203_),
    .A1(_1899_),
    .A2(net606));
 sg13g2_nand2_1 _3088_ (.Y(_1199_),
    .A(net98),
    .B(_1193_));
 sg13g2_o21ai_1 _3089_ (.B1(_1199_),
    .Y(_0204_),
    .A1(_1898_),
    .A2(net607));
 sg13g2_nand2_1 _3090_ (.Y(_1200_),
    .A(net139),
    .B(net607));
 sg13g2_o21ai_1 _3091_ (.B1(_1200_),
    .Y(_0205_),
    .A1(_1901_),
    .A2(net607));
 sg13g2_nand2_1 _3092_ (.Y(_1201_),
    .A(net141),
    .B(net607));
 sg13g2_o21ai_1 _3093_ (.B1(_1201_),
    .Y(_0206_),
    .A1(net717),
    .A2(net607));
 sg13g2_nand4_1 _3094_ (.B(net822),
    .C(net820),
    .A(net737),
    .Y(_1202_),
    .D(_1134_));
 sg13g2_nand2_1 _3095_ (.Y(_1203_),
    .A(net78),
    .B(_1202_));
 sg13g2_o21ai_1 _3096_ (.B1(_1203_),
    .Y(_0207_),
    .A1(net708),
    .A2(_1151_));
 sg13g2_nand2_1 _3097_ (.Y(_1204_),
    .A(net246),
    .B(_1202_));
 sg13g2_o21ai_1 _3098_ (.B1(_1204_),
    .Y(_0208_),
    .A1(net708),
    .A2(_1153_));
 sg13g2_nand2_1 _3099_ (.Y(_1205_),
    .A(net132),
    .B(_1202_));
 sg13g2_o21ai_1 _3100_ (.B1(_1205_),
    .Y(_0209_),
    .A1(net708),
    .A2(_1155_));
 sg13g2_nand2_1 _3101_ (.Y(_1206_),
    .A(net195),
    .B(_1202_));
 sg13g2_o21ai_1 _3102_ (.B1(_1206_),
    .Y(_0210_),
    .A1(net708),
    .A2(_1157_));
 sg13g2_nand2_1 _3103_ (.Y(_1207_),
    .A(net64),
    .B(_1202_));
 sg13g2_o21ai_1 _3104_ (.B1(_1207_),
    .Y(_0211_),
    .A1(net708),
    .A2(_1159_));
 sg13g2_nand2_1 _3105_ (.Y(_1208_),
    .A(net108),
    .B(_1202_));
 sg13g2_o21ai_1 _3106_ (.B1(_1208_),
    .Y(_0212_),
    .A1(net709),
    .A2(_1161_));
 sg13g2_nand2_1 _3107_ (.Y(_1209_),
    .A(net197),
    .B(_1202_));
 sg13g2_o21ai_1 _3108_ (.B1(_1209_),
    .Y(_0213_),
    .A1(net708),
    .A2(_1163_));
 sg13g2_nand2_1 _3109_ (.Y(_1210_),
    .A(net112),
    .B(_1202_));
 sg13g2_o21ai_1 _3110_ (.B1(_1210_),
    .Y(_0214_),
    .A1(net709),
    .A2(_1165_));
 sg13g2_and4_1 _3111_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .B(net820),
    .C(_1964_),
    .D(_1136_),
    .X(_1211_));
 sg13g2_nor2_1 _3112_ (.A(net362),
    .B(net604),
    .Y(_1212_));
 sg13g2_a21oi_1 _3113_ (.A1(_1168_),
    .A2(net604),
    .Y(_0215_),
    .B1(_1212_));
 sg13g2_nor2_1 _3114_ (.A(net416),
    .B(net604),
    .Y(_1213_));
 sg13g2_a21oi_1 _3115_ (.A1(_1170_),
    .A2(net604),
    .Y(_0216_),
    .B1(_1213_));
 sg13g2_nor2_1 _3116_ (.A(net276),
    .B(net604),
    .Y(_1214_));
 sg13g2_a21oi_1 _3117_ (.A1(_1172_),
    .A2(net604),
    .Y(_0217_),
    .B1(_1214_));
 sg13g2_nor2_1 _3118_ (.A(net325),
    .B(net604),
    .Y(_1215_));
 sg13g2_a21oi_1 _3119_ (.A1(_1173_),
    .A2(net604),
    .Y(_0218_),
    .B1(_1215_));
 sg13g2_nor2_1 _3120_ (.A(net323),
    .B(net605),
    .Y(_1216_));
 sg13g2_a21oi_1 _3121_ (.A1(_1176_),
    .A2(net605),
    .Y(_0219_),
    .B1(_1216_));
 sg13g2_nor2_1 _3122_ (.A(net499),
    .B(_1211_),
    .Y(_1217_));
 sg13g2_a21oi_1 _3123_ (.A1(_1178_),
    .A2(net605),
    .Y(_0220_),
    .B1(net500));
 sg13g2_nor2_1 _3124_ (.A(net329),
    .B(net605),
    .Y(_1218_));
 sg13g2_a21oi_1 _3125_ (.A1(_1180_),
    .A2(net605),
    .Y(_0221_),
    .B1(_1218_));
 sg13g2_nor2_1 _3126_ (.A(net272),
    .B(net605),
    .Y(_1219_));
 sg13g2_a21oi_1 _3127_ (.A1(_1182_),
    .A2(net605),
    .Y(_0222_),
    .B1(_1219_));
 sg13g2_nand4_1 _3128_ (.B(net820),
    .C(_1964_),
    .A(net737),
    .Y(_1220_),
    .D(_1183_));
 sg13g2_nand2_1 _3129_ (.Y(_1221_),
    .A(net223),
    .B(net627));
 sg13g2_o21ai_1 _3130_ (.B1(_1221_),
    .Y(_0223_),
    .A1(net721),
    .A2(net627));
 sg13g2_nand2_1 _3131_ (.Y(_1222_),
    .A(net199),
    .B(net627));
 sg13g2_o21ai_1 _3132_ (.B1(_1222_),
    .Y(_0224_),
    .A1(net720),
    .A2(net627));
 sg13g2_nand2_1 _3133_ (.Y(_1223_),
    .A(net175),
    .B(net627));
 sg13g2_o21ai_1 _3134_ (.B1(_1223_),
    .Y(_0225_),
    .A1(net718),
    .A2(net627));
 sg13g2_nand2_1 _3135_ (.Y(_1224_),
    .A(net164),
    .B(net629));
 sg13g2_o21ai_1 _3136_ (.B1(_1224_),
    .Y(_0226_),
    .A1(net719),
    .A2(net629));
 sg13g2_nand2_1 _3137_ (.Y(_1225_),
    .A(net248),
    .B(net627));
 sg13g2_o21ai_1 _3138_ (.B1(_1225_),
    .Y(_0227_),
    .A1(_1899_),
    .A2(net627));
 sg13g2_nand2_1 _3139_ (.Y(_1226_),
    .A(net167),
    .B(net628));
 sg13g2_o21ai_1 _3140_ (.B1(_1226_),
    .Y(_0228_),
    .A1(_1898_),
    .A2(net628));
 sg13g2_nand2_1 _3141_ (.Y(_1227_),
    .A(net128),
    .B(net629));
 sg13g2_o21ai_1 _3142_ (.B1(_1227_),
    .Y(_0229_),
    .A1(_1901_),
    .A2(net629));
 sg13g2_nand2_1 _3143_ (.Y(_1228_),
    .A(net161),
    .B(net628));
 sg13g2_o21ai_1 _3144_ (.B1(_1228_),
    .Y(_0230_),
    .A1(net717),
    .A2(net628));
 sg13g2_nand2_2 _3145_ (.Y(_1229_),
    .A(net735),
    .B(_1148_));
 sg13g2_nand3_1 _3146_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .C(_1148_),
    .A(net735),
    .Y(_1230_));
 sg13g2_nand2_1 _3147_ (.Y(_1231_),
    .A(net118),
    .B(_1230_));
 sg13g2_o21ai_1 _3148_ (.B1(_1231_),
    .Y(_0231_),
    .A1(_1168_),
    .A2(_1229_));
 sg13g2_nand2_1 _3149_ (.Y(_1232_),
    .A(net145),
    .B(_1230_));
 sg13g2_o21ai_1 _3150_ (.B1(_1232_),
    .Y(_0232_),
    .A1(_1170_),
    .A2(_1229_));
 sg13g2_nand2_1 _3151_ (.Y(_1233_),
    .A(net120),
    .B(_1230_));
 sg13g2_o21ai_1 _3152_ (.B1(_1233_),
    .Y(_0233_),
    .A1(_1172_),
    .A2(_1229_));
 sg13g2_nand2_1 _3153_ (.Y(_1234_),
    .A(net193),
    .B(_1230_));
 sg13g2_o21ai_1 _3154_ (.B1(_1234_),
    .Y(_0234_),
    .A1(_1173_),
    .A2(_1229_));
 sg13g2_nand2_1 _3155_ (.Y(_1235_),
    .A(net100),
    .B(_1230_));
 sg13g2_o21ai_1 _3156_ (.B1(_1235_),
    .Y(_0235_),
    .A1(_1176_),
    .A2(_1229_));
 sg13g2_nand2_1 _3157_ (.Y(_1236_),
    .A(net134),
    .B(_1230_));
 sg13g2_o21ai_1 _3158_ (.B1(_1236_),
    .Y(_0236_),
    .A1(_1178_),
    .A2(_1229_));
 sg13g2_nand2_1 _3159_ (.Y(_1237_),
    .A(net116),
    .B(_1230_));
 sg13g2_o21ai_1 _3160_ (.B1(_1237_),
    .Y(_0237_),
    .A1(_1180_),
    .A2(_1229_));
 sg13g2_nand2_1 _3161_ (.Y(_1238_),
    .A(net143),
    .B(_1230_));
 sg13g2_o21ai_1 _3162_ (.B1(_1238_),
    .Y(_0238_),
    .A1(_1182_),
    .A2(_1229_));
 sg13g2_nand3_1 _3163_ (.B(net633),
    .C(_0609_),
    .A(net739),
    .Y(_1239_));
 sg13g2_a21oi_1 _3164_ (.A1(net1070),
    .A2(_1148_),
    .Y(_1240_),
    .B1(net822));
 sg13g2_xor2_1 _3165_ (.B(_1240_),
    .A(net814),
    .X(_1241_));
 sg13g2_xor2_1 _3166_ (.B(net1015),
    .A(net822),
    .X(_1242_));
 sg13g2_nand3_1 _3167_ (.B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .C(_1183_),
    .A(net820),
    .Y(_1243_));
 sg13g2_xnor2_1 _3168_ (.Y(_1244_),
    .A(net810),
    .B(_1242_));
 sg13g2_xnor2_1 _3169_ (.Y(_1245_),
    .A(net708),
    .B(_1183_));
 sg13g2_xnor2_1 _3170_ (.Y(_1246_),
    .A(net807),
    .B(_1245_));
 sg13g2_nand3_1 _3171_ (.B(_1244_),
    .C(_1246_),
    .A(_1243_),
    .Y(_1247_));
 sg13g2_a21oi_1 _3172_ (.A1(net820),
    .A2(_1183_),
    .Y(_1248_),
    .B1(net1017));
 sg13g2_nand2b_1 _3173_ (.Y(_1249_),
    .B(_1243_),
    .A_N(_1148_));
 sg13g2_nor2_1 _3174_ (.A(_1248_),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_xor2_1 _3175_ (.B(_1250_),
    .A(net806),
    .X(_1251_));
 sg13g2_nor3_1 _3176_ (.A(_1241_),
    .B(_1247_),
    .C(_1251_),
    .Y(_1252_));
 sg13g2_o21ai_1 _3177_ (.B1(_0735_),
    .Y(_1253_),
    .A1(net768),
    .A2(_1252_));
 sg13g2_nand2b_1 _3178_ (.Y(_1254_),
    .B(_1253_),
    .A_N(_1239_));
 sg13g2_nand2_1 _3179_ (.Y(_1255_),
    .A(_0735_),
    .B(_1240_));
 sg13g2_mux2_1 _3180_ (.A0(net822),
    .A1(net955),
    .S(net768),
    .X(_1256_));
 sg13g2_a22oi_1 _3181_ (.Y(_1257_),
    .B1(_0606_),
    .B2(_1256_),
    .A2(net955),
    .A1(net749));
 sg13g2_a21oi_1 _3182_ (.A1(_1255_),
    .A2(_1257_),
    .Y(_1258_),
    .B1(net578));
 sg13g2_a21o_1 _3183_ (.A2(net578),
    .A1(net822),
    .B1(_1258_),
    .X(_0239_));
 sg13g2_nand2_1 _3184_ (.Y(_1259_),
    .A(net768),
    .B(net968));
 sg13g2_o21ai_1 _3185_ (.B1(_1259_),
    .Y(_1260_),
    .A1(net768),
    .A2(_1962_));
 sg13g2_nand2_1 _3186_ (.Y(_1261_),
    .A(_0735_),
    .B(_1242_));
 sg13g2_a22oi_1 _3187_ (.Y(_1262_),
    .B1(_0606_),
    .B2(_1260_),
    .A2(net968),
    .A1(net749));
 sg13g2_a21oi_1 _3188_ (.A1(_1261_),
    .A2(_1262_),
    .Y(_1263_),
    .B1(net578));
 sg13g2_a21o_1 _3189_ (.A2(net578),
    .A1(net1015),
    .B1(_1263_),
    .X(_0240_));
 sg13g2_nand2_1 _3190_ (.Y(_1264_),
    .A(net768),
    .B(net983));
 sg13g2_o21ai_1 _3191_ (.B1(_1264_),
    .Y(_1265_),
    .A1(net768),
    .A2(net709));
 sg13g2_nand2_1 _3192_ (.Y(_1266_),
    .A(_0735_),
    .B(_1245_));
 sg13g2_a22oi_1 _3193_ (.Y(_1267_),
    .B1(_0606_),
    .B2(_1265_),
    .A2(net983),
    .A1(net749));
 sg13g2_a21oi_1 _3194_ (.A1(_1266_),
    .A2(_1267_),
    .Y(_1268_),
    .B1(net578));
 sg13g2_a21o_1 _3195_ (.A2(_1254_),
    .A1(net820),
    .B1(_1268_),
    .X(_0241_));
 sg13g2_nand2_1 _3196_ (.Y(_1269_),
    .A(_0735_),
    .B(_1250_));
 sg13g2_nand2_1 _3197_ (.Y(_1270_),
    .A(net768),
    .B(net960));
 sg13g2_o21ai_1 _3198_ (.B1(_1270_),
    .Y(_1271_),
    .A1(net768),
    .A2(_1964_));
 sg13g2_a22oi_1 _3199_ (.Y(_1272_),
    .B1(_0606_),
    .B2(_1271_),
    .A2(net960),
    .A1(net749));
 sg13g2_a21oi_1 _3200_ (.A1(_1269_),
    .A2(_1272_),
    .Y(_1273_),
    .B1(net578));
 sg13g2_a21o_1 _3201_ (.A2(net578),
    .A1(net1017),
    .B1(_1273_),
    .X(_0242_));
 sg13g2_nor2b_2 _3202_ (.A(_0966_),
    .B_N(_0967_),
    .Y(_1274_));
 sg13g2_nand2b_1 _3203_ (.Y(_1275_),
    .B(_0967_),
    .A_N(_0966_));
 sg13g2_nor2_1 _3204_ (.A(net404),
    .B(_1274_),
    .Y(_1276_));
 sg13g2_mux4_1 _3205_ (.S0(net815),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .S1(net811),
    .X(_1277_));
 sg13g2_nand2b_2 _3206_ (.Y(_1278_),
    .B(net811),
    .A_N(net808));
 sg13g2_nor2_2 _3207_ (.A(net809),
    .B(net807),
    .Y(_1279_));
 sg13g2_mux2_1 _3208_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .S(net815),
    .X(_1280_));
 sg13g2_nor2_1 _3209_ (.A(net815),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .Y(_1281_));
 sg13g2_nor2b_1 _3210_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .B_N(net815),
    .Y(_1282_));
 sg13g2_nor3_1 _3211_ (.A(_1278_),
    .B(_1281_),
    .C(_1282_),
    .Y(_1283_));
 sg13g2_a221oi_1 _3212_ (.B2(_1280_),
    .C1(_1283_),
    .B1(_1279_),
    .A1(net808),
    .Y(_1284_),
    .A2(_1277_));
 sg13g2_nor2_1 _3213_ (.A(net805),
    .B(_1284_),
    .Y(_1285_));
 sg13g2_nand2_1 _3214_ (.Y(_1286_),
    .A(net806),
    .B(_1279_));
 sg13g2_nor2_1 _3215_ (.A(net812),
    .B(_1286_),
    .Y(_1287_));
 sg13g2_a21oi_1 _3216_ (.A1(net118),
    .A2(_1287_),
    .Y(_1288_),
    .B1(_1285_));
 sg13g2_a21oi_1 _3217_ (.A1(_1274_),
    .A2(_1288_),
    .Y(_0243_),
    .B1(net405));
 sg13g2_mux4_1 _3218_ (.S0(net815),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .S1(net811),
    .X(_1289_));
 sg13g2_mux2_1 _3219_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .S(net816),
    .X(_1290_));
 sg13g2_nor2b_1 _3220_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .B_N(net815),
    .Y(_1291_));
 sg13g2_nor2_1 _3221_ (.A(net815),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ),
    .Y(_1292_));
 sg13g2_nor3_1 _3222_ (.A(_1278_),
    .B(_1291_),
    .C(_1292_),
    .Y(_1293_));
 sg13g2_a221oi_1 _3223_ (.B2(_1279_),
    .C1(_1293_),
    .B1(_1290_),
    .A1(net808),
    .Y(_1294_),
    .A2(_1289_));
 sg13g2_nor3_1 _3224_ (.A(net805),
    .B(net601),
    .C(_1294_),
    .Y(_1295_));
 sg13g2_and2_1 _3225_ (.A(_1274_),
    .B(_1287_),
    .X(_1296_));
 sg13g2_a22oi_1 _3226_ (.Y(_1297_),
    .B1(_1296_),
    .B2(net145),
    .A2(net601),
    .A1(net894));
 sg13g2_nand2b_1 _3227_ (.Y(_0244_),
    .B(_1297_),
    .A_N(_1295_));
 sg13g2_mux4_1 _3228_ (.S0(net817),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .S1(net811),
    .X(_1298_));
 sg13g2_nor2_1 _3229_ (.A(net817),
    .B(net321),
    .Y(_1299_));
 sg13g2_nor2b_1 _3230_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[26] ),
    .B_N(net815),
    .Y(_1300_));
 sg13g2_nor3_1 _3231_ (.A(_1278_),
    .B(_1299_),
    .C(_1300_),
    .Y(_1301_));
 sg13g2_mux2_1 _3232_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .S(net817),
    .X(_1302_));
 sg13g2_a221oi_1 _3233_ (.B2(_1279_),
    .C1(_1301_),
    .B1(_1302_),
    .A1(net808),
    .Y(_1303_),
    .A2(_1298_));
 sg13g2_nor3_1 _3234_ (.A(net805),
    .B(net601),
    .C(_1303_),
    .Y(_1304_));
 sg13g2_a22oi_1 _3235_ (.Y(_1305_),
    .B1(_1296_),
    .B2(net120),
    .A2(net601),
    .A1(net495));
 sg13g2_nand2b_1 _3236_ (.Y(_0245_),
    .B(_1305_),
    .A_N(_1304_));
 sg13g2_mux2_1 _3237_ (.A0(net325),
    .A1(net164),
    .S(net812),
    .X(_1306_));
 sg13g2_nand2b_1 _3238_ (.Y(_1307_),
    .B(net812),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ));
 sg13g2_o21ai_1 _3239_ (.B1(_1307_),
    .Y(_1308_),
    .A1(net812),
    .A2(net77));
 sg13g2_or2_1 _3240_ (.X(_1309_),
    .B(net63),
    .A(net812));
 sg13g2_o21ai_1 _3241_ (.B1(net807),
    .Y(_1310_),
    .A1(net809),
    .A2(_1308_));
 sg13g2_a21oi_1 _3242_ (.A1(net809),
    .A2(_1306_),
    .Y(_1311_),
    .B1(_1310_));
 sg13g2_mux2_1 _3243_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .S(net812),
    .X(_1312_));
 sg13g2_a21oi_1 _3244_ (.A1(net813),
    .A2(_1978_),
    .Y(_1313_),
    .B1(net809));
 sg13g2_a221oi_1 _3245_ (.B2(_1309_),
    .C1(net807),
    .B1(_1313_),
    .A1(net809),
    .Y(_1314_),
    .A2(_1312_));
 sg13g2_nor4_1 _3246_ (.A(net806),
    .B(net601),
    .C(_1311_),
    .D(_1314_),
    .Y(_1315_));
 sg13g2_a22oi_1 _3247_ (.Y(_1316_),
    .B1(_1296_),
    .B2(net193),
    .A2(net601),
    .A1(net559));
 sg13g2_nand2b_1 _3248_ (.Y(_0246_),
    .B(_1316_),
    .A_N(_1315_));
 sg13g2_mux4_1 _3249_ (.S0(net816),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .S1(net811),
    .X(_1317_));
 sg13g2_mux2_1 _3250_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .S(net816),
    .X(_1318_));
 sg13g2_nor2b_1 _3251_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[28] ),
    .B_N(net816),
    .Y(_1319_));
 sg13g2_nor2_1 _3252_ (.A(net816),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .Y(_1320_));
 sg13g2_nor3_1 _3253_ (.A(_1278_),
    .B(_1319_),
    .C(_1320_),
    .Y(_1321_));
 sg13g2_a221oi_1 _3254_ (.B2(_1279_),
    .C1(_1321_),
    .B1(_1318_),
    .A1(net808),
    .Y(_1322_),
    .A2(_1317_));
 sg13g2_nor3_1 _3255_ (.A(net805),
    .B(net601),
    .C(_1322_),
    .Y(_1323_));
 sg13g2_a22oi_1 _3256_ (.Y(_1324_),
    .B1(_1296_),
    .B2(net100),
    .A2(net601),
    .A1(net544));
 sg13g2_nand2b_1 _3257_ (.Y(_0247_),
    .B(_1324_),
    .A_N(_1323_));
 sg13g2_mux4_1 _3258_ (.S0(net818),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .S1(net811),
    .X(_1325_));
 sg13g2_nor2_1 _3259_ (.A(net818),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .Y(_1326_));
 sg13g2_nor2b_1 _3260_ (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[29] ),
    .B_N(net818),
    .Y(_1327_));
 sg13g2_nor3_1 _3261_ (.A(_1278_),
    .B(_1326_),
    .C(_1327_),
    .Y(_1328_));
 sg13g2_mux2_1 _3262_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .S(net818),
    .X(_1329_));
 sg13g2_a221oi_1 _3263_ (.B2(_1279_),
    .C1(_1328_),
    .B1(_1329_),
    .A1(net808),
    .Y(_1330_),
    .A2(_1325_));
 sg13g2_nor3_1 _3264_ (.A(net805),
    .B(net602),
    .C(_1330_),
    .Y(_1331_));
 sg13g2_a22oi_1 _3265_ (.Y(_1332_),
    .B1(_1296_),
    .B2(net134),
    .A2(net602),
    .A1(net897));
 sg13g2_nand2b_1 _3266_ (.Y(_0248_),
    .B(_1332_),
    .A_N(_1331_));
 sg13g2_nand2b_1 _3267_ (.Y(_1333_),
    .B(net814),
    .A_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ));
 sg13g2_o21ai_1 _3268_ (.B1(_1333_),
    .Y(_1334_),
    .A1(net814),
    .A2(net139));
 sg13g2_mux2_1 _3269_ (.A0(net329),
    .A1(net128),
    .S(net814),
    .X(_1335_));
 sg13g2_or2_1 _3270_ (.X(_1336_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[6] ),
    .A(net813));
 sg13g2_o21ai_1 _3271_ (.B1(net807),
    .Y(_1337_),
    .A1(net810),
    .A2(_1334_));
 sg13g2_a21oi_1 _3272_ (.A1(net809),
    .A2(_1335_),
    .Y(_1338_),
    .B1(_1337_));
 sg13g2_mux2_1 _3273_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .S(net813),
    .X(_1339_));
 sg13g2_a21oi_1 _3274_ (.A1(net813),
    .A2(_1979_),
    .Y(_1340_),
    .B1(net809));
 sg13g2_a221oi_1 _3275_ (.B2(_1336_),
    .C1(net807),
    .B1(_1340_),
    .A1(net810),
    .Y(_1341_),
    .A2(_1339_));
 sg13g2_nor4_1 _3276_ (.A(net805),
    .B(net602),
    .C(_1338_),
    .D(_1341_),
    .Y(_1342_));
 sg13g2_a22oi_1 _3277_ (.Y(_1343_),
    .B1(_1296_),
    .B2(net116),
    .A2(net602),
    .A1(net876));
 sg13g2_nand2b_1 _3278_ (.Y(_0249_),
    .B(_1343_),
    .A_N(_1342_));
 sg13g2_mux4_1 _3279_ (.S0(net818),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .S1(net811),
    .X(_1344_));
 sg13g2_nor2_1 _3280_ (.A(net819),
    .B(net314),
    .Y(_1345_));
 sg13g2_nor2b_1 _3281_ (.A(net201),
    .B_N(net818),
    .Y(_1346_));
 sg13g2_nor3_1 _3282_ (.A(_1278_),
    .B(_1345_),
    .C(_1346_),
    .Y(_1347_));
 sg13g2_mux2_1 _3283_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .S(net818),
    .X(_1348_));
 sg13g2_a221oi_1 _3284_ (.B2(_1279_),
    .C1(_1347_),
    .B1(_1348_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .Y(_1349_),
    .A2(_1344_));
 sg13g2_nor3_1 _3285_ (.A(net805),
    .B(net602),
    .C(_1349_),
    .Y(_1350_));
 sg13g2_a22oi_1 _3286_ (.Y(_1351_),
    .B1(_1296_),
    .B2(net143),
    .A2(net602),
    .A1(net874));
 sg13g2_nand2b_1 _3287_ (.Y(_0250_),
    .B(_1351_),
    .A_N(_1350_));
 sg13g2_nor3_2 _3288_ (.A(net749),
    .B(_0605_),
    .C(_1239_),
    .Y(_1352_));
 sg13g2_mux2_1 _3289_ (.A0(net955),
    .A1(_1256_),
    .S(_1352_),
    .X(_0251_));
 sg13g2_mux2_1 _3290_ (.A0(net968),
    .A1(_1260_),
    .S(_1352_),
    .X(_0252_));
 sg13g2_mux2_1 _3291_ (.A0(net983),
    .A1(_1265_),
    .S(_1352_),
    .X(_0253_));
 sg13g2_mux2_1 _3292_ (.A0(net960),
    .A1(_1271_),
    .S(_1352_),
    .X(_0254_));
 sg13g2_a21oi_1 _3293_ (.A1(_1274_),
    .A2(_1286_),
    .Y(_1353_),
    .B1(net812));
 sg13g2_a21oi_1 _3294_ (.A1(net814),
    .A2(_1274_),
    .Y(_0255_),
    .B1(_1353_));
 sg13g2_nand3_1 _3295_ (.B(net810),
    .C(_1274_),
    .A(net819),
    .Y(_1354_));
 sg13g2_a21o_1 _3296_ (.A2(_1274_),
    .A1(net819),
    .B1(net810),
    .X(_1355_));
 sg13g2_and2_1 _3297_ (.A(_1354_),
    .B(_1355_),
    .X(_0256_));
 sg13g2_nand4_1 _3298_ (.B(net809),
    .C(net807),
    .A(net812),
    .Y(_1356_),
    .D(_1274_));
 sg13g2_xnor2_1 _3299_ (.Y(_0257_),
    .A(net808),
    .B(_1354_));
 sg13g2_xor2_1 _3300_ (.B(_1356_),
    .A(net805),
    .X(_1357_));
 sg13g2_nor2_1 _3301_ (.A(_1296_),
    .B(_1357_),
    .Y(_0258_));
 sg13g2_nand2_2 _3302_ (.Y(_1358_),
    .A(_1123_),
    .B(_1129_));
 sg13g2_nand3_1 _3303_ (.B(net301),
    .C(net631),
    .A(net1046),
    .Y(_1359_));
 sg13g2_nor4_1 _3304_ (.A(net803),
    .B(net794),
    .C(net790),
    .D(_1914_),
    .Y(_1360_));
 sg13g2_a21o_1 _3305_ (.A2(net631),
    .A1(\u_usb_cdc.sie_in_req ),
    .B1(net626),
    .X(_1361_));
 sg13g2_o21ai_1 _3306_ (.B1(_1359_),
    .Y(_1362_),
    .A1(net803),
    .A2(_1361_));
 sg13g2_nor2_1 _3307_ (.A(_1358_),
    .B(_1362_),
    .Y(_1363_));
 sg13g2_a21oi_1 _3308_ (.A1(_1912_),
    .A2(_1358_),
    .Y(_0259_),
    .B1(_1363_));
 sg13g2_xnor2_1 _3309_ (.Y(_1364_),
    .A(net803),
    .B(net795));
 sg13g2_nand2_1 _3310_ (.Y(_1365_),
    .A(_1128_),
    .B(_1364_));
 sg13g2_o21ai_1 _3311_ (.B1(_1365_),
    .Y(_1366_),
    .A1(net927),
    .A2(_1128_));
 sg13g2_nand2_1 _3312_ (.Y(_1367_),
    .A(net795),
    .B(_1358_));
 sg13g2_o21ai_1 _3313_ (.B1(net1027),
    .Y(_0260_),
    .A1(_1358_),
    .A2(_1366_));
 sg13g2_nand3_1 _3314_ (.B(net795),
    .C(net790),
    .A(net803),
    .Y(_1368_));
 sg13g2_a21o_1 _3315_ (.A2(net795),
    .A1(net803),
    .B1(net790),
    .X(_1369_));
 sg13g2_and2_1 _3316_ (.A(_1368_),
    .B(_1369_),
    .X(_1370_));
 sg13g2_mux2_1 _3317_ (.A0(net280),
    .A1(_1370_),
    .S(_1128_),
    .X(_1371_));
 sg13g2_nor2_1 _3318_ (.A(_1358_),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_a21oi_1 _3319_ (.A1(_1913_),
    .A2(_1358_),
    .Y(_0261_),
    .B1(_1372_));
 sg13g2_nand3_1 _3320_ (.B(net335),
    .C(net632),
    .A(net1046),
    .Y(_1373_));
 sg13g2_xnor2_1 _3321_ (.Y(_1374_),
    .A(_1914_),
    .B(_1368_));
 sg13g2_o21ai_1 _3322_ (.B1(_1373_),
    .Y(_1375_),
    .A1(_1361_),
    .A2(_1374_));
 sg13g2_mux2_1 _3323_ (.A0(_1375_),
    .A1(net788),
    .S(_1358_),
    .X(_0262_));
 sg13g2_nor2_1 _3324_ (.A(net619),
    .B(_0662_),
    .Y(_1376_));
 sg13g2_nor2_2 _3325_ (.A(_0724_),
    .B(_1376_),
    .Y(_1377_));
 sg13g2_nor2_1 _3326_ (.A(net518),
    .B(net569),
    .Y(_1378_));
 sg13g2_a21oi_1 _3327_ (.A1(_1894_),
    .A2(net569),
    .Y(_0263_),
    .B1(_1378_));
 sg13g2_nor2_1 _3328_ (.A(net423),
    .B(net569),
    .Y(_1379_));
 sg13g2_a21oi_1 _3329_ (.A1(net720),
    .A2(_1377_),
    .Y(_0264_),
    .B1(_1379_));
 sg13g2_nor2_1 _3330_ (.A(net341),
    .B(net569),
    .Y(_1380_));
 sg13g2_a21oi_1 _3331_ (.A1(net718),
    .A2(net569),
    .Y(_0265_),
    .B1(_1380_));
 sg13g2_nor2_1 _3332_ (.A(net271),
    .B(net569),
    .Y(_1381_));
 sg13g2_a21oi_1 _3333_ (.A1(net719),
    .A2(net569),
    .Y(_0266_),
    .B1(_1381_));
 sg13g2_nor2_1 _3334_ (.A(net479),
    .B(_1377_),
    .Y(_1382_));
 sg13g2_a21oi_1 _3335_ (.A1(net717),
    .A2(net569),
    .Y(_0267_),
    .B1(_1382_));
 sg13g2_nor2b_1 _3336_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .B_N(net841),
    .Y(_1383_));
 sg13g2_nor3_2 _3337_ (.A(_0614_),
    .B(_0639_),
    .C(_1383_),
    .Y(_1384_));
 sg13g2_nand2_1 _3338_ (.Y(_1385_),
    .A(net269),
    .B(_1384_));
 sg13g2_o21ai_1 _3339_ (.B1(_1385_),
    .Y(_0268_),
    .A1(_1954_),
    .A2(_1384_));
 sg13g2_mux2_1 _3340_ (.A0(net880),
    .A1(net391),
    .S(_1384_),
    .X(_0269_));
 sg13g2_mux2_1 _3341_ (.A0(net926),
    .A1(net392),
    .S(_1384_),
    .X(_0270_));
 sg13g2_mux2_1 _3342_ (.A0(net905),
    .A1(net510),
    .S(_1384_),
    .X(_0271_));
 sg13g2_mux2_1 _3343_ (.A0(net896),
    .A1(net384),
    .S(_1384_),
    .X(_0272_));
 sg13g2_mux2_1 _3344_ (.A0(net865),
    .A1(net458),
    .S(_1384_),
    .X(_0273_));
 sg13g2_mux2_1 _3345_ (.A0(net886),
    .A1(net364),
    .S(_1384_),
    .X(_0274_));
 sg13g2_nand2_1 _3346_ (.Y(_1386_),
    .A(net738),
    .B(net619));
 sg13g2_o21ai_1 _3347_ (.B1(_1386_),
    .Y(_1387_),
    .A1(net751),
    .A2(_0778_));
 sg13g2_and2_1 _3348_ (.A(_0723_),
    .B(_1387_),
    .X(_1388_));
 sg13g2_nor2_1 _3349_ (.A(net269),
    .B(net570),
    .Y(_1389_));
 sg13g2_a21oi_1 _3350_ (.A1(_1894_),
    .A2(net570),
    .Y(_0275_),
    .B1(_1389_));
 sg13g2_nor2_1 _3351_ (.A(net391),
    .B(net570),
    .Y(_1390_));
 sg13g2_a21oi_1 _3352_ (.A1(_1895_),
    .A2(net570),
    .Y(_0276_),
    .B1(_1390_));
 sg13g2_nor2_1 _3353_ (.A(net392),
    .B(net570),
    .Y(_1391_));
 sg13g2_a21oi_1 _3354_ (.A1(net718),
    .A2(net571),
    .Y(_0277_),
    .B1(_1391_));
 sg13g2_nor2_1 _3355_ (.A(net510),
    .B(net570),
    .Y(_1392_));
 sg13g2_a21oi_1 _3356_ (.A1(net719),
    .A2(net570),
    .Y(_0278_),
    .B1(_1392_));
 sg13g2_nor2_1 _3357_ (.A(net384),
    .B(net570),
    .Y(_1393_));
 sg13g2_a21oi_1 _3358_ (.A1(_1899_),
    .A2(net571),
    .Y(_0279_),
    .B1(_1393_));
 sg13g2_nor2_1 _3359_ (.A(net458),
    .B(net571),
    .Y(_1394_));
 sg13g2_a21oi_1 _3360_ (.A1(_1898_),
    .A2(net571),
    .Y(_0280_),
    .B1(_1394_));
 sg13g2_nor2_1 _3361_ (.A(net364),
    .B(net571),
    .Y(_1395_));
 sg13g2_a21oi_1 _3362_ (.A1(_1901_),
    .A2(net571),
    .Y(_0281_),
    .B1(_1395_));
 sg13g2_o21ai_1 _3363_ (.B1(_1386_),
    .Y(_1396_),
    .A1(_0710_),
    .A2(_0784_));
 sg13g2_and2_1 _3364_ (.A(_0723_),
    .B(_1396_),
    .X(_1397_));
 sg13g2_mux2_1 _3365_ (.A0(net415),
    .A1(_0711_),
    .S(_1397_),
    .X(_0282_));
 sg13g2_or2_1 _3366_ (.X(_0283_),
    .B(_1397_),
    .A(net345));
 sg13g2_a21oi_1 _3367_ (.A1(_0653_),
    .A2(_0705_),
    .Y(_1398_),
    .B1(net620));
 sg13g2_nor2_2 _3368_ (.A(_0724_),
    .B(_1398_),
    .Y(_1399_));
 sg13g2_nor2_1 _3369_ (.A(net920),
    .B(_1399_),
    .Y(_1400_));
 sg13g2_a21oi_1 _3370_ (.A1(net721),
    .A2(_1399_),
    .Y(_0284_),
    .B1(_1400_));
 sg13g2_nor2_1 _3371_ (.A(net910),
    .B(_1399_),
    .Y(_1401_));
 sg13g2_a21oi_1 _3372_ (.A1(net720),
    .A2(_1399_),
    .Y(_0285_),
    .B1(_1401_));
 sg13g2_nor2_1 _3373_ (.A(net884),
    .B(_1399_),
    .Y(_1402_));
 sg13g2_a21oi_1 _3374_ (.A1(_1898_),
    .A2(_1399_),
    .Y(_0286_),
    .B1(_1402_));
 sg13g2_nor2_1 _3375_ (.A(net993),
    .B(_1399_),
    .Y(_1403_));
 sg13g2_a21oi_1 _3376_ (.A1(_1900_),
    .A2(_1399_),
    .Y(_0287_),
    .B1(_1403_));
 sg13g2_nor3_1 _3377_ (.A(_0673_),
    .B(net617),
    .C(_0752_),
    .Y(_1404_));
 sg13g2_nor3_1 _3378_ (.A(net620),
    .B(_0675_),
    .C(_1404_),
    .Y(_1405_));
 sg13g2_nor2_1 _3379_ (.A(_0724_),
    .B(_1405_),
    .Y(_1406_));
 sg13g2_nor2_1 _3380_ (.A(net864),
    .B(net568),
    .Y(_1407_));
 sg13g2_o21ai_1 _3381_ (.B1(_0673_),
    .Y(_1408_),
    .A1(_1900_),
    .A2(_0752_));
 sg13g2_nor2_1 _3382_ (.A(net761),
    .B(_1408_),
    .Y(_1409_));
 sg13g2_a21oi_1 _3383_ (.A1(net567),
    .A2(_1409_),
    .Y(_0288_),
    .B1(_1407_));
 sg13g2_nor2_1 _3384_ (.A(net856),
    .B(net567),
    .Y(_1410_));
 sg13g2_nor2_1 _3385_ (.A(net757),
    .B(_1408_),
    .Y(_1411_));
 sg13g2_a21oi_1 _3386_ (.A1(net567),
    .A2(_1411_),
    .Y(_0289_),
    .B1(_1410_));
 sg13g2_nor2_1 _3387_ (.A(net523),
    .B(net567),
    .Y(_1412_));
 sg13g2_nor2_1 _3388_ (.A(net756),
    .B(_1408_),
    .Y(_1413_));
 sg13g2_a21oi_1 _3389_ (.A1(net567),
    .A2(_1413_),
    .Y(_0290_),
    .B1(_1412_));
 sg13g2_nor2_1 _3390_ (.A(net916),
    .B(net567),
    .Y(_1414_));
 sg13g2_nor2_1 _3391_ (.A(net755),
    .B(_1408_),
    .Y(_1415_));
 sg13g2_a21oi_1 _3392_ (.A1(net568),
    .A2(_1415_),
    .Y(_0291_),
    .B1(_1414_));
 sg13g2_nor2_1 _3393_ (.A(net538),
    .B(net567),
    .Y(_1416_));
 sg13g2_nor2_1 _3394_ (.A(net754),
    .B(_1408_),
    .Y(_1417_));
 sg13g2_a21oi_1 _3395_ (.A1(net568),
    .A2(_1417_),
    .Y(_0292_),
    .B1(_1416_));
 sg13g2_nor2_1 _3396_ (.A(net854),
    .B(net567),
    .Y(_1418_));
 sg13g2_nor2_1 _3397_ (.A(net753),
    .B(_1408_),
    .Y(_1419_));
 sg13g2_a21oi_1 _3398_ (.A1(net568),
    .A2(_1419_),
    .Y(_0293_),
    .B1(_1418_));
 sg13g2_nor2_1 _3399_ (.A(net890),
    .B(net568),
    .Y(_1420_));
 sg13g2_nor2_1 _3400_ (.A(\u_usb_cdc.sie_out_data[6] ),
    .B(_1408_),
    .Y(_1421_));
 sg13g2_a21oi_1 _3401_ (.A1(net568),
    .A2(_1421_),
    .Y(_0294_),
    .B1(_1420_));
 sg13g2_a21oi_1 _3402_ (.A1(_0554_),
    .A2(_0640_),
    .Y(_1422_),
    .B1(_1920_));
 sg13g2_nor2_1 _3403_ (.A(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .B(_1422_),
    .Y(_1423_));
 sg13g2_o21ai_1 _3404_ (.B1(_0647_),
    .Y(_1424_),
    .A1(_0844_),
    .A2(_1423_));
 sg13g2_a21oi_1 _3405_ (.A1(_0558_),
    .A2(_0605_),
    .Y(_1425_),
    .B1(\u_usb_cdc.u_ctrl_endp.state_q[6] ));
 sg13g2_or3_1 _3406_ (.A(_0844_),
    .B(_1424_),
    .C(_1425_),
    .X(_1426_));
 sg13g2_nor2_1 _3407_ (.A(_1915_),
    .B(_1424_),
    .Y(_1427_));
 sg13g2_a21oi_1 _3408_ (.A1(_1915_),
    .A2(_1426_),
    .Y(_0295_),
    .B1(_1427_));
 sg13g2_nand2_1 _3409_ (.Y(_1428_),
    .A(net785),
    .B(_1424_));
 sg13g2_nor2_1 _3410_ (.A(_0548_),
    .B(_0660_),
    .Y(_1429_));
 sg13g2_nand2_1 _3411_ (.Y(_1430_),
    .A(_0549_),
    .B(_0661_));
 sg13g2_o21ai_1 _3412_ (.B1(_1428_),
    .Y(_0296_),
    .A1(_1426_),
    .A2(_1430_));
 sg13g2_nand2_1 _3413_ (.Y(_1431_),
    .A(net783),
    .B(_1424_));
 sg13g2_xor2_1 _3414_ (.B(_0549_),
    .A(net783),
    .X(_1432_));
 sg13g2_o21ai_1 _3415_ (.B1(_1431_),
    .Y(_0297_),
    .A1(_1426_),
    .A2(_1432_));
 sg13g2_nand2_1 _3416_ (.Y(_1433_),
    .A(net778),
    .B(_1424_));
 sg13g2_nand3_1 _3417_ (.B(net778),
    .C(_0548_),
    .A(net783),
    .Y(_1434_));
 sg13g2_nand3b_1 _3418_ (.B(_1434_),
    .C(_0665_),
    .Y(_1435_),
    .A_N(_1426_));
 sg13g2_nand2_1 _3419_ (.Y(_0298_),
    .A(_1433_),
    .B(_1435_));
 sg13g2_nand2_1 _3420_ (.Y(_1436_),
    .A(net775),
    .B(_1424_));
 sg13g2_nand4_1 _3421_ (.B(net778),
    .C(net775),
    .A(net783),
    .Y(_1437_),
    .D(_0548_));
 sg13g2_xor2_1 _3422_ (.B(_1434_),
    .A(net775),
    .X(_1438_));
 sg13g2_o21ai_1 _3423_ (.B1(_1436_),
    .Y(_0299_),
    .A1(_1426_),
    .A2(_1438_));
 sg13g2_nand2_1 _3424_ (.Y(_1439_),
    .A(net772),
    .B(_1424_));
 sg13g2_nand2_1 _3425_ (.Y(_1440_),
    .A(net775),
    .B(net772));
 sg13g2_nor2_1 _3426_ (.A(_1434_),
    .B(_1440_),
    .Y(_1441_));
 sg13g2_xor2_1 _3427_ (.B(_1437_),
    .A(net772),
    .X(_1442_));
 sg13g2_o21ai_1 _3428_ (.B1(_1439_),
    .Y(_0300_),
    .A1(_1426_),
    .A2(_1442_));
 sg13g2_nand2_1 _3429_ (.Y(_1443_),
    .A(net951),
    .B(_1424_));
 sg13g2_xnor2_1 _3430_ (.Y(_1444_),
    .A(net951),
    .B(_1441_));
 sg13g2_o21ai_1 _3431_ (.B1(_1443_),
    .Y(_0301_),
    .A1(_1426_),
    .A2(_1444_));
 sg13g2_nand2b_1 _3432_ (.Y(_1445_),
    .B(_1239_),
    .A_N(net769));
 sg13g2_and2_1 _3433_ (.A(net578),
    .B(_1445_),
    .X(_0302_));
 sg13g2_nor2_1 _3434_ (.A(net942),
    .B(_0869_),
    .Y(_1446_));
 sg13g2_a21oi_1 _3435_ (.A1(_1906_),
    .A2(net582),
    .Y(_0303_),
    .B1(_1446_));
 sg13g2_nor2_1 _3436_ (.A(net766),
    .B(net582),
    .Y(_1447_));
 sg13g2_a21oi_1 _3437_ (.A1(_1907_),
    .A2(net582),
    .Y(_0304_),
    .B1(_1447_));
 sg13g2_mux2_1 _3438_ (.A0(net764),
    .A1(net1002),
    .S(net582),
    .X(_0305_));
 sg13g2_nor2_1 _3439_ (.A(net762),
    .B(net582),
    .Y(_1448_));
 sg13g2_a21oi_1 _3440_ (.A1(_1908_),
    .A2(_0869_),
    .Y(_0306_),
    .B1(_1448_));
 sg13g2_nand2_1 _3441_ (.Y(_1449_),
    .A(net252),
    .B(net580));
 sg13g2_o21ai_1 _3442_ (.B1(_1449_),
    .Y(_0307_),
    .A1(_1895_),
    .A2(net580));
 sg13g2_nand2_1 _3443_ (.Y(_1450_),
    .A(net213),
    .B(net580));
 sg13g2_o21ai_1 _3444_ (.B1(_1450_),
    .Y(_0308_),
    .A1(net718),
    .A2(net581));
 sg13g2_nand2_1 _3445_ (.Y(_1451_),
    .A(net200),
    .B(net580));
 sg13g2_o21ai_1 _3446_ (.B1(_1451_),
    .Y(_0309_),
    .A1(net719),
    .A2(net580));
 sg13g2_nand2_1 _3447_ (.Y(_1452_),
    .A(net237),
    .B(net581));
 sg13g2_o21ai_1 _3448_ (.B1(_1452_),
    .Y(_0310_),
    .A1(_1899_),
    .A2(net581));
 sg13g2_nand2_1 _3449_ (.Y(_1453_),
    .A(net214),
    .B(net580));
 sg13g2_o21ai_1 _3450_ (.B1(_1453_),
    .Y(_0311_),
    .A1(_1898_),
    .A2(net581));
 sg13g2_nand2_1 _3451_ (.Y(_1454_),
    .A(net250),
    .B(net580));
 sg13g2_o21ai_1 _3452_ (.B1(_1454_),
    .Y(_0312_),
    .A1(_1901_),
    .A2(net580));
 sg13g2_a21oi_1 _3453_ (.A1(_1932_),
    .A2(_1383_),
    .Y(_1455_),
    .B1(_0614_));
 sg13g2_a22oi_1 _3454_ (.Y(_1456_),
    .B1(_0647_),
    .B2(_1455_),
    .A2(net878),
    .A1(net738));
 sg13g2_nor4_1 _3455_ (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[2] ),
    .B(\u_usb_cdc.u_ctrl_endp.addr_dd[5] ),
    .C(\u_usb_cdc.u_ctrl_endp.addr_dd[4] ),
    .D(\u_usb_cdc.u_ctrl_endp.addr_dd[6] ),
    .Y(_1457_));
 sg13g2_nor4_1 _3456_ (.A(\u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .B(\u_usb_cdc.u_ctrl_endp.addr_dd[1] ),
    .C(\u_usb_cdc.u_ctrl_endp.addr_dd[0] ),
    .D(\u_usb_cdc.u_ctrl_endp.addr_dd[3] ),
    .Y(_1458_));
 sg13g2_a21oi_1 _3457_ (.A1(_1457_),
    .A2(_1458_),
    .Y(_1459_),
    .B1(net878));
 sg13g2_o21ai_1 _3458_ (.B1(_1459_),
    .Y(_1460_),
    .A1(net415),
    .A2(_1932_));
 sg13g2_mux2_1 _3459_ (.A0(_1460_),
    .A1(net937),
    .S(_1456_),
    .X(_0313_));
 sg13g2_nand2_1 _3460_ (.Y(_1461_),
    .A(net346),
    .B(_1456_));
 sg13g2_o21ai_1 _3461_ (.B1(_1459_),
    .Y(_1462_),
    .A1(_1932_),
    .A2(net345));
 sg13g2_o21ai_1 _3462_ (.B1(net347),
    .Y(_0314_),
    .A1(_1456_),
    .A2(_1462_));
 sg13g2_nor2b_1 _3463_ (.A(net739),
    .B_N(net1046),
    .Y(_1463_));
 sg13g2_nor3_1 _3464_ (.A(_0589_),
    .B(_0591_),
    .C(_0976_),
    .Y(_1464_));
 sg13g2_a21o_1 _3465_ (.A2(_1464_),
    .A1(_0494_),
    .B1(_1463_),
    .X(_0315_));
 sg13g2_nor3_2 _3466_ (.A(net833),
    .B(net832),
    .C(net837),
    .Y(_1465_));
 sg13g2_nand4_1 _3467_ (.B(net507),
    .C(net1005),
    .A(net460),
    .Y(_1466_),
    .D(_1465_));
 sg13g2_nand3_1 _3468_ (.B(net742),
    .C(_1466_),
    .A(net1005),
    .Y(_1467_));
 sg13g2_nor2_1 _3469_ (.A(net712),
    .B(_1465_),
    .Y(_1468_));
 sg13g2_o21ai_1 _3470_ (.B1(_1467_),
    .Y(_1469_),
    .A1(net1005),
    .A2(net742));
 sg13g2_nor2_1 _3471_ (.A(_1468_),
    .B(_1469_),
    .Y(_0316_));
 sg13g2_a21oi_1 _3472_ (.A1(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .A2(net742),
    .Y(_1470_),
    .B1(net507));
 sg13g2_nand3_1 _3473_ (.B(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .C(net742),
    .A(net507),
    .Y(_1471_));
 sg13g2_nor2_1 _3474_ (.A(net460),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_nor3_1 _3475_ (.A(_1468_),
    .B(net508),
    .C(_1472_),
    .Y(_0317_));
 sg13g2_a21oi_1 _3476_ (.A1(_1921_),
    .A2(_1471_),
    .Y(_0318_),
    .B1(_1468_));
 sg13g2_nand2_1 _3477_ (.Y(_1473_),
    .A(net289),
    .B(net594));
 sg13g2_o21ai_1 _3478_ (.B1(_1473_),
    .Y(_0319_),
    .A1(net289),
    .A2(_0894_));
 sg13g2_nand2_1 _3479_ (.Y(_1474_),
    .A(net319),
    .B(net594));
 sg13g2_xnor2_1 _3480_ (.Y(_1475_),
    .A(net319),
    .B(net289));
 sg13g2_o21ai_1 _3481_ (.B1(_1474_),
    .Y(_0320_),
    .A1(_0894_),
    .A2(_1475_));
 sg13g2_nand2_1 _3482_ (.Y(_1476_),
    .A(net230),
    .B(net594));
 sg13g2_a21o_1 _3483_ (.A2(\u_usb_cdc.u_sie.in_byte_q[0] ),
    .A1(\u_usb_cdc.u_sie.in_byte_q[1] ),
    .B1(net230),
    .X(_1477_));
 sg13g2_nand2_1 _3484_ (.Y(_1478_),
    .A(_0611_),
    .B(_1477_));
 sg13g2_o21ai_1 _3485_ (.B1(_1476_),
    .Y(_0321_),
    .A1(_0894_),
    .A2(_1478_));
 sg13g2_nand2_1 _3486_ (.Y(_1479_),
    .A(net339),
    .B(net594));
 sg13g2_xor2_1 _3487_ (.B(_0611_),
    .A(net339),
    .X(_1480_));
 sg13g2_o21ai_1 _3488_ (.B1(_1479_),
    .Y(_0322_),
    .A1(_0894_),
    .A2(_1480_));
 sg13g2_nor2_1 _3489_ (.A(net835),
    .B(net839),
    .Y(_1481_));
 sg13g2_nor3_1 _3490_ (.A(net834),
    .B(net839),
    .C(net836),
    .Y(_1482_));
 sg13g2_a21o_1 _3491_ (.A2(_1482_),
    .A1(_0905_),
    .B1(_0595_),
    .X(_1483_));
 sg13g2_nor3_2 _3492_ (.A(net840),
    .B(net836),
    .C(net577),
    .Y(_1484_));
 sg13g2_xor2_1 _3493_ (.B(_0514_),
    .A(_0500_),
    .X(_1485_));
 sg13g2_a22oi_1 _3494_ (.Y(_0323_),
    .B1(net573),
    .B2(_1485_),
    .A2(net576),
    .A1(_1946_));
 sg13g2_a22oi_1 _3495_ (.Y(_0324_),
    .B1(net573),
    .B2(_0514_),
    .A2(net576),
    .A1(_1947_));
 sg13g2_a22oi_1 _3496_ (.Y(_0325_),
    .B1(net572),
    .B2(_0520_),
    .A2(net575),
    .A1(_1949_));
 sg13g2_a22oi_1 _3497_ (.Y(_0326_),
    .B1(net572),
    .B2(_0503_),
    .A2(net575),
    .A1(_1948_));
 sg13g2_a22oi_1 _3498_ (.Y(_0327_),
    .B1(net572),
    .B2(net445),
    .A2(net575),
    .A1(_1951_));
 sg13g2_a22oi_1 _3499_ (.Y(_0328_),
    .B1(net572),
    .B2(net549),
    .A2(net575),
    .A1(_1950_));
 sg13g2_a22oi_1 _3500_ (.Y(_0329_),
    .B1(net573),
    .B2(_0506_),
    .A2(net576),
    .A1(_1953_));
 sg13g2_a22oi_1 _3501_ (.Y(_0330_),
    .B1(_1484_),
    .B2(_0521_),
    .A2(net576),
    .A1(_1952_));
 sg13g2_a22oi_1 _3502_ (.Y(_0331_),
    .B1(net573),
    .B2(_0516_),
    .A2(net577),
    .A1(_1945_));
 sg13g2_a22oi_1 _3503_ (.Y(_0332_),
    .B1(net572),
    .B2(_0517_),
    .A2(net575),
    .A1(_1944_));
 sg13g2_a22oi_1 _3504_ (.Y(_0333_),
    .B1(net573),
    .B2(_1949_),
    .A2(net575),
    .A1(_1943_));
 sg13g2_a22oi_1 _3505_ (.Y(_0334_),
    .B1(net572),
    .B2(_1948_),
    .A2(net577),
    .A1(_1942_));
 sg13g2_a22oi_1 _3506_ (.Y(_0335_),
    .B1(net572),
    .B2(_1951_),
    .A2(net575),
    .A1(_1941_));
 sg13g2_a22oi_1 _3507_ (.Y(_0336_),
    .B1(net572),
    .B2(_1950_),
    .A2(net575),
    .A1(_1940_));
 sg13g2_a22oi_1 _3508_ (.Y(_0337_),
    .B1(net573),
    .B2(_1953_),
    .A2(net576),
    .A1(_1939_));
 sg13g2_xnor2_1 _3509_ (.Y(_1486_),
    .A(_1952_),
    .B(_1485_));
 sg13g2_a22oi_1 _3510_ (.Y(_0338_),
    .B1(net573),
    .B2(_1486_),
    .A2(net576),
    .A1(_1938_));
 sg13g2_nand2_1 _3511_ (.Y(_1487_),
    .A(net766),
    .B(net594));
 sg13g2_nor2_1 _3512_ (.A(net747),
    .B(_1481_),
    .Y(_1488_));
 sg13g2_or2_1 _3513_ (.X(_1489_),
    .B(_1481_),
    .A(net747));
 sg13g2_nor2b_1 _3514_ (.A(net799),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .Y(_1490_));
 sg13g2_a21oi_1 _3515_ (.A1(net799),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .Y(_1491_),
    .B1(_1490_));
 sg13g2_mux2_1 _3516_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .S(net797),
    .X(_1492_));
 sg13g2_a21oi_1 _3517_ (.A1(net792),
    .A2(_1492_),
    .Y(_1493_),
    .B1(net789));
 sg13g2_o21ai_1 _3518_ (.B1(_1493_),
    .Y(_1494_),
    .A1(net792),
    .A2(_1491_));
 sg13g2_a21oi_1 _3519_ (.A1(net799),
    .A2(_1967_),
    .Y(_1495_),
    .B1(net792));
 sg13g2_o21ai_1 _3520_ (.B1(_1495_),
    .Y(_1496_),
    .A1(net799),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ));
 sg13g2_mux2_1 _3521_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .S(net797),
    .X(_1497_));
 sg13g2_a21oi_1 _3522_ (.A1(net792),
    .A2(_1497_),
    .Y(_1498_),
    .B1(_1913_));
 sg13g2_a21oi_1 _3523_ (.A1(_1496_),
    .A2(_1498_),
    .Y(_1499_),
    .B1(net788));
 sg13g2_a22oi_1 _3524_ (.Y(_1500_),
    .B1(_1494_),
    .B2(_1499_),
    .A2(net626),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ));
 sg13g2_o21ai_1 _3525_ (.B1(net625),
    .Y(_1501_),
    .A1(_0576_),
    .A2(_1500_));
 sg13g2_nor2b_1 _3526_ (.A(net773),
    .B_N(net770),
    .Y(_1502_));
 sg13g2_nand2b_1 _3527_ (.Y(_1503_),
    .B(net770),
    .A_N(net773));
 sg13g2_nand2_1 _3528_ (.Y(_1504_),
    .A(net780),
    .B(_0651_));
 sg13g2_a21oi_1 _3529_ (.A1(net780),
    .A2(_0651_),
    .Y(_1505_),
    .B1(net776));
 sg13g2_nor2_1 _3530_ (.A(_0664_),
    .B(_1505_),
    .Y(_1506_));
 sg13g2_nand2b_1 _3531_ (.Y(_1507_),
    .B(_1429_),
    .A_N(net780));
 sg13g2_nand2b_1 _3532_ (.Y(_1508_),
    .B(_1507_),
    .A_N(_0551_));
 sg13g2_o21ai_1 _3533_ (.B1(_1502_),
    .Y(_1509_),
    .A1(_1506_),
    .A2(_1508_));
 sg13g2_and2_1 _3534_ (.A(net777),
    .B(_0547_),
    .X(_1510_));
 sg13g2_nand2_1 _3535_ (.Y(_1511_),
    .A(net716),
    .B(net782));
 sg13g2_a21oi_1 _3536_ (.A1(_0547_),
    .A2(_1511_),
    .Y(_1512_),
    .B1(net777));
 sg13g2_o21ai_1 _3537_ (.B1(_0544_),
    .Y(_1513_),
    .A1(_1510_),
    .A2(_1512_));
 sg13g2_nand3_1 _3538_ (.B(net777),
    .C(_0549_),
    .A(net780),
    .Y(_1514_));
 sg13g2_a21oi_1 _3539_ (.A1(_0650_),
    .A2(_0661_),
    .Y(_1515_),
    .B1(_1440_));
 sg13g2_nand2_2 _3540_ (.Y(_1516_),
    .A(_1917_),
    .B(\u_usb_cdc.u_ctrl_endp.req_q[8] ));
 sg13g2_inv_1 _3541_ (.Y(_1517_),
    .A(_1516_));
 sg13g2_a21oi_1 _3542_ (.A1(_1514_),
    .A2(_1515_),
    .Y(_1518_),
    .B1(_1516_));
 sg13g2_nor3_2 _3543_ (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .B(net779),
    .C(_0547_),
    .Y(_1519_));
 sg13g2_a21oi_1 _3544_ (.A1(net787),
    .A2(net716),
    .Y(_1520_),
    .B1(_0543_));
 sg13g2_o21ai_1 _3545_ (.B1(_0552_),
    .Y(_1521_),
    .A1(_1519_),
    .A2(_1520_));
 sg13g2_nand4_1 _3546_ (.B(_1513_),
    .C(_1518_),
    .A(_1509_),
    .Y(_1522_),
    .D(_1521_));
 sg13g2_a22oi_1 _3547_ (.Y(_1523_),
    .B1(_1519_),
    .B2(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .A2(\u_usb_cdc.configured_o ),
    .A1(\u_usb_cdc.u_ctrl_endp.req_q[4] ));
 sg13g2_nand3_1 _3548_ (.B(_1504_),
    .C(_1507_),
    .A(net776),
    .Y(_1524_));
 sg13g2_nor2_1 _3549_ (.A(net774),
    .B(_1918_),
    .Y(_1525_));
 sg13g2_nand2b_1 _3550_ (.Y(_1526_),
    .B(_1525_),
    .A_N(_1524_));
 sg13g2_nand3_1 _3551_ (.B(_1523_),
    .C(_1526_),
    .A(_1522_),
    .Y(_1527_));
 sg13g2_and3_2 _3552_ (.X(_1528_),
    .A(_0554_),
    .B(_0560_),
    .C(_0576_));
 sg13g2_nand3_1 _3553_ (.B(_0560_),
    .C(_0576_),
    .A(_0554_),
    .Y(_1529_));
 sg13g2_a21oi_1 _3554_ (.A1(_1527_),
    .A2(_1528_),
    .Y(_1530_),
    .B1(_1501_));
 sg13g2_o21ai_1 _3555_ (.B1(net597),
    .Y(_1531_),
    .A1(net967),
    .A2(net624));
 sg13g2_o21ai_1 _3556_ (.B1(_1487_),
    .Y(_0339_),
    .A1(_1530_),
    .A2(_1531_));
 sg13g2_nand2_1 _3557_ (.Y(_1532_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .B(net626));
 sg13g2_mux4_1 _3558_ (.S0(net797),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .S1(net792),
    .X(_1533_));
 sg13g2_a21oi_1 _3559_ (.A1(net799),
    .A2(_1968_),
    .Y(_1534_),
    .B1(net792));
 sg13g2_o21ai_1 _3560_ (.B1(_1534_),
    .Y(_1535_),
    .A1(net797),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ));
 sg13g2_mux2_1 _3561_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .S(net797),
    .X(_1536_));
 sg13g2_a21oi_1 _3562_ (.A1(net792),
    .A2(_1536_),
    .Y(_1537_),
    .B1(_1913_));
 sg13g2_nand2_1 _3563_ (.Y(_1538_),
    .A(_1535_),
    .B(_1537_));
 sg13g2_o21ai_1 _3564_ (.B1(_1538_),
    .Y(_1539_),
    .A1(net789),
    .A2(_1533_));
 sg13g2_o21ai_1 _3565_ (.B1(_1532_),
    .Y(_1540_),
    .A1(net788),
    .A2(_1539_));
 sg13g2_a21oi_1 _3566_ (.A1(net631),
    .A2(_1540_),
    .Y(_1541_),
    .B1(_1489_));
 sg13g2_nor2b_1 _3567_ (.A(_0660_),
    .B_N(net781),
    .Y(_1542_));
 sg13g2_o21ai_1 _3568_ (.B1(net778),
    .Y(_1543_),
    .A1(_0705_),
    .A2(_1542_));
 sg13g2_or2_1 _3569_ (.X(_1544_),
    .B(_0705_),
    .A(net776));
 sg13g2_or2_1 _3570_ (.X(_1545_),
    .B(_1544_),
    .A(_1542_));
 sg13g2_o21ai_1 _3571_ (.B1(_1504_),
    .Y(_1546_),
    .A1(net780),
    .A2(_0548_));
 sg13g2_a21oi_1 _3572_ (.A1(_1543_),
    .A2(_1545_),
    .Y(_1547_),
    .B1(_0668_));
 sg13g2_a21oi_1 _3573_ (.A1(_1546_),
    .A2(_1547_),
    .Y(_1548_),
    .B1(net770));
 sg13g2_o21ai_1 _3574_ (.B1(net776),
    .Y(_1549_),
    .A1(net781),
    .A2(_1429_));
 sg13g2_nand3b_1 _3575_ (.B(_0542_),
    .C(_0664_),
    .Y(_1550_),
    .A_N(net776));
 sg13g2_a21oi_1 _3576_ (.A1(_1549_),
    .A2(_1550_),
    .Y(_1551_),
    .B1(_1503_));
 sg13g2_a221oi_1 _3577_ (.B2(_1430_),
    .C1(_1440_),
    .B1(_1510_),
    .A1(_0541_),
    .Y(_1552_),
    .A2(_1505_));
 sg13g2_nor4_1 _3578_ (.A(_1516_),
    .B(_1548_),
    .C(_1551_),
    .D(_1552_),
    .Y(_1553_));
 sg13g2_nor3_1 _3579_ (.A(net777),
    .B(_0550_),
    .C(_0660_),
    .Y(_1554_));
 sg13g2_nor4_1 _3580_ (.A(net774),
    .B(_1918_),
    .C(_1510_),
    .D(_1554_),
    .Y(_1555_));
 sg13g2_o21ai_1 _3581_ (.B1(_1528_),
    .Y(_1556_),
    .A1(_1553_),
    .A2(_1555_));
 sg13g2_o21ai_1 _3582_ (.B1(net597),
    .Y(_1557_),
    .A1(net940),
    .A2(net624));
 sg13g2_a21oi_1 _3583_ (.A1(_1541_),
    .A2(_1556_),
    .Y(_1558_),
    .B1(_1557_));
 sg13g2_a21o_1 _3584_ (.A2(net594),
    .A1(net765),
    .B1(_1558_),
    .X(_0340_));
 sg13g2_nand2_1 _3585_ (.Y(_1559_),
    .A(net763),
    .B(net594));
 sg13g2_nand2_1 _3586_ (.Y(_1560_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .B(net626));
 sg13g2_mux4_1 _3587_ (.S0(net798),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .S1(net791),
    .X(_1561_));
 sg13g2_a21oi_1 _3588_ (.A1(net800),
    .A2(_1969_),
    .Y(_1562_),
    .B1(net791));
 sg13g2_o21ai_1 _3589_ (.B1(_1562_),
    .Y(_1563_),
    .A1(net798),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ));
 sg13g2_mux2_1 _3590_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .S(net798),
    .X(_1564_));
 sg13g2_a21oi_1 _3591_ (.A1(net791),
    .A2(_1564_),
    .Y(_1565_),
    .B1(_1913_));
 sg13g2_nand2_1 _3592_ (.Y(_1566_),
    .A(_1563_),
    .B(_1565_));
 sg13g2_o21ai_1 _3593_ (.B1(_1566_),
    .Y(_1567_),
    .A1(net789),
    .A2(_1561_));
 sg13g2_o21ai_1 _3594_ (.B1(_1560_),
    .Y(_1568_),
    .A1(net788),
    .A2(_1567_));
 sg13g2_a21oi_1 _3595_ (.A1(_0541_),
    .A2(_0549_),
    .Y(_1569_),
    .B1(net776));
 sg13g2_a21oi_1 _3596_ (.A1(net716),
    .A2(_1510_),
    .Y(_1570_),
    .B1(_1569_));
 sg13g2_a21oi_1 _3597_ (.A1(net776),
    .A2(_1546_),
    .Y(_1571_),
    .B1(_0551_));
 sg13g2_nor2b_1 _3598_ (.A(_1570_),
    .B_N(net774),
    .Y(_1572_));
 sg13g2_nor2_1 _3599_ (.A(_0542_),
    .B(_0670_),
    .Y(_1573_));
 sg13g2_nor3_1 _3600_ (.A(net771),
    .B(_1572_),
    .C(_1573_),
    .Y(_1574_));
 sg13g2_a21oi_1 _3601_ (.A1(net773),
    .A2(_1511_),
    .Y(_1575_),
    .B1(_0650_));
 sg13g2_a21oi_1 _3602_ (.A1(_0650_),
    .A2(_1429_),
    .Y(_1576_),
    .B1(_1575_));
 sg13g2_a21oi_1 _3603_ (.A1(net770),
    .A2(_1576_),
    .Y(_1577_),
    .B1(_1516_));
 sg13g2_o21ai_1 _3604_ (.B1(_1577_),
    .Y(_1578_),
    .A1(_1503_),
    .A2(_1571_));
 sg13g2_nor2_1 _3605_ (.A(_1574_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_a221oi_1 _3606_ (.B2(_1528_),
    .C1(_1489_),
    .B1(_1579_),
    .A1(net631),
    .Y(_1580_),
    .A2(_1568_));
 sg13g2_o21ai_1 _3607_ (.B1(net597),
    .Y(_1581_),
    .A1(net945),
    .A2(net624));
 sg13g2_o21ai_1 _3608_ (.B1(_1559_),
    .Y(_0341_),
    .A1(_1580_),
    .A2(_1581_));
 sg13g2_nand2_1 _3609_ (.Y(_1582_),
    .A(net1011),
    .B(net593));
 sg13g2_nand2_1 _3610_ (.Y(_1583_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .B(net626));
 sg13g2_mux4_1 _3611_ (.S0(net797),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .S1(net791),
    .X(_1584_));
 sg13g2_a21oi_1 _3612_ (.A1(net800),
    .A2(_1970_),
    .Y(_1585_),
    .B1(net791));
 sg13g2_o21ai_1 _3613_ (.B1(_1585_),
    .Y(_1586_),
    .A1(net800),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ));
 sg13g2_mux2_1 _3614_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .S(net798),
    .X(_1587_));
 sg13g2_a21oi_1 _3615_ (.A1(net791),
    .A2(_1587_),
    .Y(_1588_),
    .B1(_1913_));
 sg13g2_nand2_1 _3616_ (.Y(_1589_),
    .A(_1586_),
    .B(_1588_));
 sg13g2_o21ai_1 _3617_ (.B1(_1589_),
    .Y(_1590_),
    .A1(net789),
    .A2(_1584_));
 sg13g2_o21ai_1 _3618_ (.B1(_1583_),
    .Y(_1591_),
    .A1(net788),
    .A2(_1590_));
 sg13g2_nand3_1 _3619_ (.B(_1525_),
    .C(_1549_),
    .A(_0665_),
    .Y(_1592_));
 sg13g2_nor2_1 _3620_ (.A(net773),
    .B(_0669_),
    .Y(_1593_));
 sg13g2_a21oi_1 _3621_ (.A1(_0547_),
    .A2(_1511_),
    .Y(_1594_),
    .B1(_1917_));
 sg13g2_nor2b_1 _3622_ (.A(_0544_),
    .B_N(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .Y(_1595_));
 sg13g2_o21ai_1 _3623_ (.B1(_1595_),
    .Y(_1596_),
    .A1(_0738_),
    .A2(_1593_));
 sg13g2_or2_1 _3624_ (.X(_1597_),
    .B(_1596_),
    .A(_1594_));
 sg13g2_o21ai_1 _3625_ (.B1(net778),
    .Y(_1598_),
    .A1(net786),
    .A2(net781));
 sg13g2_o21ai_1 _3626_ (.B1(_1502_),
    .Y(_1599_),
    .A1(_1542_),
    .A2(_1598_));
 sg13g2_o21ai_1 _3627_ (.B1(_1599_),
    .Y(_1600_),
    .A1(net771),
    .A2(_1544_));
 sg13g2_o21ai_1 _3628_ (.B1(_1592_),
    .Y(_1601_),
    .A1(_1597_),
    .A2(_1600_));
 sg13g2_a221oi_1 _3629_ (.B2(_1528_),
    .C1(_1489_),
    .B1(_1601_),
    .A1(net631),
    .Y(_1602_),
    .A2(_1591_));
 sg13g2_o21ai_1 _3630_ (.B1(net597),
    .Y(_1603_),
    .A1(net966),
    .A2(net624));
 sg13g2_o21ai_1 _3631_ (.B1(_1582_),
    .Y(_0342_),
    .A1(_1602_),
    .A2(_1603_));
 sg13g2_nand2_1 _3632_ (.Y(_1604_),
    .A(net980),
    .B(net593));
 sg13g2_nor2b_1 _3633_ (.A(net800),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .Y(_1605_));
 sg13g2_a21oi_1 _3634_ (.A1(net799),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .Y(_1606_),
    .B1(_1605_));
 sg13g2_mux2_1 _3635_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .S(net801),
    .X(_1607_));
 sg13g2_a21oi_1 _3636_ (.A1(net796),
    .A2(_1607_),
    .Y(_1608_),
    .B1(net790));
 sg13g2_o21ai_1 _3637_ (.B1(_1608_),
    .Y(_1609_),
    .A1(net793),
    .A2(_1606_));
 sg13g2_a21oi_1 _3638_ (.A1(net799),
    .A2(_1971_),
    .Y(_1610_),
    .B1(net793));
 sg13g2_o21ai_1 _3639_ (.B1(_1610_),
    .Y(_1611_),
    .A1(net799),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ));
 sg13g2_mux2_1 _3640_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .S(net801),
    .X(_1612_));
 sg13g2_a21oi_1 _3641_ (.A1(net793),
    .A2(_1612_),
    .Y(_1613_),
    .B1(_1913_));
 sg13g2_a21oi_1 _3642_ (.A1(_1611_),
    .A2(_1613_),
    .Y(_1614_),
    .B1(net788));
 sg13g2_a22oi_1 _3643_ (.Y(_1615_),
    .B1(_1609_),
    .B2(_1614_),
    .A2(net626),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ));
 sg13g2_nor3_1 _3644_ (.A(net781),
    .B(_0549_),
    .C(_0670_),
    .Y(_1616_));
 sg13g2_nor2b_1 _3645_ (.A(_1616_),
    .B_N(net771),
    .Y(_1617_));
 sg13g2_nor2_1 _3646_ (.A(_1516_),
    .B(_1617_),
    .Y(_1618_));
 sg13g2_a22oi_1 _3647_ (.Y(_1619_),
    .B1(_0850_),
    .B2(_0552_),
    .A2(_0652_),
    .A1(_0544_));
 sg13g2_and2_1 _3648_ (.A(_1525_),
    .B(_1543_),
    .X(_1620_));
 sg13g2_a22oi_1 _3649_ (.Y(_1621_),
    .B1(_1620_),
    .B2(_1544_),
    .A2(_1619_),
    .A1(_1618_));
 sg13g2_nor2_1 _3650_ (.A(_1529_),
    .B(_1621_),
    .Y(_1622_));
 sg13g2_o21ai_1 _3651_ (.B1(net625),
    .Y(_1623_),
    .A1(_0576_),
    .A2(_1615_));
 sg13g2_nor2_1 _3652_ (.A(_1622_),
    .B(_1623_),
    .Y(_1624_));
 sg13g2_o21ai_1 _3653_ (.B1(net597),
    .Y(_1625_),
    .A1(net929),
    .A2(net624));
 sg13g2_o21ai_1 _3654_ (.B1(_1604_),
    .Y(_0343_),
    .A1(_1624_),
    .A2(_1625_));
 sg13g2_nand2_1 _3655_ (.Y(_1626_),
    .A(net995),
    .B(net593));
 sg13g2_nand2_1 _3656_ (.Y(_1627_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .B(net626));
 sg13g2_mux4_1 _3657_ (.S0(net797),
    .A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .A3(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .S1(net791),
    .X(_1628_));
 sg13g2_a21oi_1 _3658_ (.A1(net800),
    .A2(_1972_),
    .Y(_1629_),
    .B1(net793));
 sg13g2_o21ai_1 _3659_ (.B1(_1629_),
    .Y(_1630_),
    .A1(net800),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ));
 sg13g2_mux2_1 _3660_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .S(net797),
    .X(_1631_));
 sg13g2_nand2_1 _3661_ (.Y(_1632_),
    .A(net791),
    .B(_1631_));
 sg13g2_nand3_1 _3662_ (.B(_1630_),
    .C(_1632_),
    .A(net789),
    .Y(_1633_));
 sg13g2_o21ai_1 _3663_ (.B1(_1633_),
    .Y(_1634_),
    .A1(net789),
    .A2(_1628_));
 sg13g2_o21ai_1 _3664_ (.B1(_1627_),
    .Y(_1635_),
    .A1(net788),
    .A2(_1634_));
 sg13g2_nor3_1 _3665_ (.A(_1918_),
    .B(_0541_),
    .C(_0670_),
    .Y(_1636_));
 sg13g2_nor2_1 _3666_ (.A(net771),
    .B(_0551_),
    .Y(_1637_));
 sg13g2_o21ai_1 _3667_ (.B1(_1637_),
    .Y(_1638_),
    .A1(_0550_),
    .A2(_1524_));
 sg13g2_nand2b_1 _3668_ (.Y(_1639_),
    .B(_1519_),
    .A_N(net773));
 sg13g2_a221oi_1 _3669_ (.B2(_1639_),
    .C1(_1516_),
    .B1(_1617_),
    .A1(_0552_),
    .Y(_1640_),
    .A2(_0850_));
 sg13g2_a22oi_1 _3670_ (.Y(_1641_),
    .B1(_1638_),
    .B2(_1640_),
    .A2(_1573_),
    .A1(\u_usb_cdc.u_ctrl_endp.req_q[2] ));
 sg13g2_a21oi_1 _3671_ (.A1(net631),
    .A2(_1635_),
    .Y(_1642_),
    .B1(_1489_));
 sg13g2_o21ai_1 _3672_ (.B1(_1642_),
    .Y(_1643_),
    .A1(_1529_),
    .A2(_1641_));
 sg13g2_o21ai_1 _3673_ (.B1(_1643_),
    .Y(_1644_),
    .A1(net992),
    .A2(net625));
 sg13g2_o21ai_1 _3674_ (.B1(_1626_),
    .Y(_0344_),
    .A1(net593),
    .A2(_1644_));
 sg13g2_nand2_1 _3675_ (.Y(_1645_),
    .A(net985),
    .B(net593));
 sg13g2_nand2_1 _3676_ (.Y(_1646_),
    .A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .B(net626));
 sg13g2_nor2b_1 _3677_ (.A(net802),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .Y(_1647_));
 sg13g2_a21oi_1 _3678_ (.A1(net802),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_mux2_1 _3679_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .S(net800),
    .X(_1649_));
 sg13g2_a21oi_1 _3680_ (.A1(net793),
    .A2(_1649_),
    .Y(_1650_),
    .B1(net789));
 sg13g2_o21ai_1 _3681_ (.B1(_1650_),
    .Y(_1651_),
    .A1(net794),
    .A2(_1648_));
 sg13g2_nor2_1 _3682_ (.A(_1912_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .Y(_1652_));
 sg13g2_nor2_1 _3683_ (.A(net802),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ),
    .Y(_1653_));
 sg13g2_nor3_1 _3684_ (.A(net794),
    .B(_1652_),
    .C(_1653_),
    .Y(_1654_));
 sg13g2_nor2_1 _3685_ (.A(_1912_),
    .B(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .Y(_1655_));
 sg13g2_o21ai_1 _3686_ (.B1(net794),
    .Y(_1656_),
    .A1(net802),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ));
 sg13g2_o21ai_1 _3687_ (.B1(net790),
    .Y(_1657_),
    .A1(_1655_),
    .A2(_1656_));
 sg13g2_o21ai_1 _3688_ (.B1(_1651_),
    .Y(_1658_),
    .A1(_1654_),
    .A2(_1657_));
 sg13g2_o21ai_1 _3689_ (.B1(_1646_),
    .Y(_1659_),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .A2(_1658_));
 sg13g2_a21oi_1 _3690_ (.A1(net785),
    .A2(_0543_),
    .Y(_1660_),
    .B1(net770));
 sg13g2_nor4_1 _3691_ (.A(_0544_),
    .B(_1516_),
    .C(_1617_),
    .D(_1660_),
    .Y(_1661_));
 sg13g2_or2_1 _3692_ (.X(_1662_),
    .B(_1661_),
    .A(_1636_));
 sg13g2_a221oi_1 _3693_ (.B2(_1528_),
    .C1(_1489_),
    .B1(_1662_),
    .A1(net631),
    .Y(_1663_),
    .A2(_1659_));
 sg13g2_o21ai_1 _3694_ (.B1(net597),
    .Y(_1664_),
    .A1(net982),
    .A2(net624));
 sg13g2_o21ai_1 _3695_ (.B1(_1645_),
    .Y(_0345_),
    .A1(_1663_),
    .A2(_1664_));
 sg13g2_nand2_1 _3696_ (.Y(_1665_),
    .A(net919),
    .B(net593));
 sg13g2_nand2_1 _3697_ (.Y(_1666_),
    .A(net491),
    .B(_1360_));
 sg13g2_a21oi_1 _3698_ (.A1(net801),
    .A2(_1973_),
    .Y(_1667_),
    .B1(net793));
 sg13g2_o21ai_1 _3699_ (.B1(_1667_),
    .Y(_1668_),
    .A1(net801),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ));
 sg13g2_mux2_1 _3700_ (.A0(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .A1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .S(net801),
    .X(_1669_));
 sg13g2_a21oi_1 _3701_ (.A1(net794),
    .A2(_1669_),
    .Y(_1670_),
    .B1(net790));
 sg13g2_nor2b_1 _3702_ (.A(net801),
    .B_N(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .Y(_1671_));
 sg13g2_a21oi_1 _3703_ (.A1(net802),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .Y(_1672_),
    .B1(_1671_));
 sg13g2_o21ai_1 _3704_ (.B1(net794),
    .Y(_1673_),
    .A1(net801),
    .A2(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ));
 sg13g2_a21oi_1 _3705_ (.A1(net801),
    .A2(_1974_),
    .Y(_1674_),
    .B1(_1673_));
 sg13g2_o21ai_1 _3706_ (.B1(net789),
    .Y(_1675_),
    .A1(net793),
    .A2(_1672_));
 sg13g2_a21oi_1 _3707_ (.A1(_1668_),
    .A2(_1670_),
    .Y(_1676_),
    .B1(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ));
 sg13g2_o21ai_1 _3708_ (.B1(_1676_),
    .Y(_1677_),
    .A1(_1674_),
    .A2(_1675_));
 sg13g2_a21oi_1 _3709_ (.A1(_1666_),
    .A2(_1677_),
    .Y(_1678_),
    .B1(_0576_));
 sg13g2_a22oi_1 _3710_ (.Y(_1679_),
    .B1(_1573_),
    .B2(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .A2(_1517_),
    .A1(_0672_));
 sg13g2_nor2_1 _3711_ (.A(_1529_),
    .B(_1679_),
    .Y(_1680_));
 sg13g2_nor3_1 _3712_ (.A(_1489_),
    .B(_1678_),
    .C(_1680_),
    .Y(_1681_));
 sg13g2_o21ai_1 _3713_ (.B1(net597),
    .Y(_1682_),
    .A1(net999),
    .A2(net624));
 sg13g2_o21ai_1 _3714_ (.B1(_1665_),
    .Y(_0346_),
    .A1(_1681_),
    .A2(_1682_));
 sg13g2_nand2_2 _3715_ (.Y(_1683_),
    .A(_1957_),
    .B(_0905_));
 sg13g2_nand3_1 _3716_ (.B(net590),
    .C(_1683_),
    .A(net766),
    .Y(_1684_));
 sg13g2_o21ai_1 _3717_ (.B1(_1684_),
    .Y(_0347_),
    .A1(_1894_),
    .A2(net598));
 sg13g2_nand3_1 _3718_ (.B(net590),
    .C(_1683_),
    .A(net764),
    .Y(_1685_));
 sg13g2_o21ai_1 _3719_ (.B1(_1685_),
    .Y(_0348_),
    .A1(_1895_),
    .A2(net598));
 sg13g2_nand3_1 _3720_ (.B(net591),
    .C(_1683_),
    .A(net762),
    .Y(_1686_));
 sg13g2_o21ai_1 _3721_ (.B1(_1686_),
    .Y(_0349_),
    .A1(_1897_),
    .A2(net598));
 sg13g2_nand3_1 _3722_ (.B(net590),
    .C(_1683_),
    .A(net1011),
    .Y(_1687_));
 sg13g2_o21ai_1 _3723_ (.B1(_1687_),
    .Y(_0350_),
    .A1(_1896_),
    .A2(net598));
 sg13g2_nand3_1 _3724_ (.B(net590),
    .C(_1683_),
    .A(net980),
    .Y(_1688_));
 sg13g2_o21ai_1 _3725_ (.B1(_1688_),
    .Y(_0351_),
    .A1(_1899_),
    .A2(net598));
 sg13g2_nand3_1 _3726_ (.B(net591),
    .C(_1683_),
    .A(net995),
    .Y(_1689_));
 sg13g2_o21ai_1 _3727_ (.B1(_1689_),
    .Y(_0352_),
    .A1(_1898_),
    .A2(net598));
 sg13g2_nand3_1 _3728_ (.B(net590),
    .C(_1683_),
    .A(net985),
    .Y(_1690_));
 sg13g2_o21ai_1 _3729_ (.B1(_1690_),
    .Y(_0353_),
    .A1(_1901_),
    .A2(net598));
 sg13g2_nand3_1 _3730_ (.B(net590),
    .C(_1683_),
    .A(net919),
    .Y(_1691_));
 sg13g2_o21ai_1 _3731_ (.B1(_1691_),
    .Y(_0354_),
    .A1(_1900_),
    .A2(net598));
 sg13g2_mux2_1 _3732_ (.A0(net761),
    .A1(net412),
    .S(net589),
    .X(_0355_));
 sg13g2_mux2_1 _3733_ (.A0(net759),
    .A1(net420),
    .S(net589),
    .X(_0356_));
 sg13g2_mux2_1 _3734_ (.A0(net756),
    .A1(net374),
    .S(net589),
    .X(_0357_));
 sg13g2_mux2_1 _3735_ (.A0(net755),
    .A1(net505),
    .S(_0602_),
    .X(_0358_));
 sg13g2_mux2_1 _3736_ (.A0(net754),
    .A1(net858),
    .S(net589),
    .X(_0359_));
 sg13g2_mux2_1 _3737_ (.A0(net753),
    .A1(net370),
    .S(net589),
    .X(_0360_));
 sg13g2_mux2_1 _3738_ (.A0(net752),
    .A1(net503),
    .S(_0602_),
    .X(_0361_));
 sg13g2_mux2_1 _3739_ (.A0(net751),
    .A1(net843),
    .S(_0602_),
    .X(_0362_));
 sg13g2_mux2_1 _3740_ (.A0(\u_usb_cdc.u_sie.data_q[0] ),
    .A1(net911),
    .S(net589),
    .X(_0363_));
 sg13g2_mux2_1 _3741_ (.A0(\u_usb_cdc.u_sie.data_q[1] ),
    .A1(net962),
    .S(net589),
    .X(_0364_));
 sg13g2_mux2_1 _3742_ (.A0(net763),
    .A1(net933),
    .S(net589),
    .X(_0365_));
 sg13g2_nor2_2 _3743_ (.A(net833),
    .B(net840),
    .Y(_1692_));
 sg13g2_inv_1 _3744_ (.Y(_1693_),
    .A(_1692_));
 sg13g2_nor2_1 _3745_ (.A(net836),
    .B(_1693_),
    .Y(_1694_));
 sg13g2_nor4_2 _3746_ (.A(_0581_),
    .B(_0599_),
    .C(_0999_),
    .Y(_1695_),
    .D(_1694_));
 sg13g2_or2_1 _3747_ (.X(_1696_),
    .B(_0618_),
    .A(_0577_));
 sg13g2_o21ai_1 _3748_ (.B1(_1696_),
    .Y(_1697_),
    .A1(_0890_),
    .A2(_1693_));
 sg13g2_mux2_1 _3749_ (.A0(net904),
    .A1(_1697_),
    .S(_1695_),
    .X(_0366_));
 sg13g2_nand2_1 _3750_ (.Y(_1698_),
    .A(_1003_),
    .B(_1692_));
 sg13g2_mux2_1 _3751_ (.A0(net957),
    .A1(_1698_),
    .S(_1695_),
    .X(_0367_));
 sg13g2_nand3_1 _3752_ (.B(_0889_),
    .C(_1692_),
    .A(net763),
    .Y(_1699_));
 sg13g2_o21ai_1 _3753_ (.B1(_1699_),
    .Y(_1700_),
    .A1(_0578_),
    .A2(_1692_));
 sg13g2_mux2_1 _3754_ (.A0(net1009),
    .A1(_1700_),
    .S(_1695_),
    .X(_0368_));
 sg13g2_o21ai_1 _3755_ (.B1(net839),
    .Y(_1701_),
    .A1(_0579_),
    .A2(_1018_));
 sg13g2_nand3_1 _3756_ (.B(_0889_),
    .C(_1692_),
    .A(net1011),
    .Y(_1702_));
 sg13g2_a22oi_1 _3757_ (.Y(_1703_),
    .B1(net633),
    .B2(net769),
    .A2(_0572_),
    .A1(\u_usb_cdc.ctrl_stall ));
 sg13g2_nand2b_1 _3758_ (.Y(_1704_),
    .B(net833),
    .A_N(_1703_));
 sg13g2_nand3_1 _3759_ (.B(_1702_),
    .C(_1704_),
    .A(_1701_),
    .Y(_1705_));
 sg13g2_mux2_1 _3760_ (.A0(net1018),
    .A1(_1705_),
    .S(_1695_),
    .X(_0369_));
 sg13g2_nor2_1 _3761_ (.A(_0529_),
    .B(_0987_),
    .Y(_1706_));
 sg13g2_nor2b_1 _3762_ (.A(_1706_),
    .B_N(_0908_),
    .Y(_1707_));
 sg13g2_nor3_1 _3763_ (.A(net748),
    .B(net750),
    .C(_1707_),
    .Y(_1708_));
 sg13g2_or2_1 _3764_ (.X(_1709_),
    .B(_1465_),
    .A(_0589_));
 sg13g2_a21oi_1 _3765_ (.A1(_1466_),
    .A2(_1709_),
    .Y(_1710_),
    .B1(net712));
 sg13g2_o21ai_1 _3766_ (.B1(_1710_),
    .Y(_1711_),
    .A1(net833),
    .A2(_1709_));
 sg13g2_nor3_1 _3767_ (.A(_1465_),
    .B(_1708_),
    .C(_1711_),
    .Y(_1712_));
 sg13g2_a21o_1 _3768_ (.A2(_1711_),
    .A1(net750),
    .B1(_1712_),
    .X(_0370_));
 sg13g2_nand2_1 _3769_ (.Y(_1713_),
    .A(_0601_),
    .B(_0623_));
 sg13g2_nor2_1 _3770_ (.A(_0466_),
    .B(_1713_),
    .Y(_1714_));
 sg13g2_a22oi_1 _3771_ (.Y(_1715_),
    .B1(_1714_),
    .B2(_0494_),
    .A2(_1706_),
    .A1(_0908_));
 sg13g2_nor4_1 _3772_ (.A(_0589_),
    .B(_0591_),
    .C(_0981_),
    .D(_1715_),
    .Y(_1716_));
 sg13g2_nor2_1 _3773_ (.A(net291),
    .B(_1716_),
    .Y(_1717_));
 sg13g2_a21oi_1 _3774_ (.A1(_1465_),
    .A2(_1710_),
    .Y(_0371_),
    .B1(net292));
 sg13g2_a22oi_1 _3775_ (.Y(_1718_),
    .B1(_0938_),
    .B2(_1936_),
    .A2(_0443_),
    .A1(net515));
 sg13g2_nor2_1 _3776_ (.A(_1937_),
    .B(_0933_),
    .Y(_1719_));
 sg13g2_nor2b_2 _3777_ (.A(_1718_),
    .B_N(_1719_),
    .Y(_1720_));
 sg13g2_a22oi_1 _3778_ (.Y(_1721_),
    .B1(_1720_),
    .B2(net531),
    .A2(net579),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ));
 sg13g2_inv_1 _3779_ (.Y(_0372_),
    .A(net532));
 sg13g2_a22oi_1 _3780_ (.Y(_1722_),
    .B1(_1720_),
    .B2(net485),
    .A2(net579),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ));
 sg13g2_inv_1 _3781_ (.Y(_0373_),
    .A(net486));
 sg13g2_a22oi_1 _3782_ (.Y(_1723_),
    .B1(_1720_),
    .B2(net899),
    .A2(net579),
    .A1(net485));
 sg13g2_inv_1 _3783_ (.Y(_0374_),
    .A(net900));
 sg13g2_a22oi_1 _3784_ (.Y(_1724_),
    .B1(_1720_),
    .B2(net527),
    .A2(net579),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ));
 sg13g2_inv_1 _3785_ (.Y(_0375_),
    .A(net528));
 sg13g2_a22oi_1 _3786_ (.Y(_1725_),
    .B1(_1720_),
    .B2(net428),
    .A2(net579),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ));
 sg13g2_inv_1 _3787_ (.Y(_0376_),
    .A(net429));
 sg13g2_a22oi_1 _3788_ (.Y(_1726_),
    .B1(_1720_),
    .B2(net862),
    .A2(_0933_),
    .A1(net428));
 sg13g2_inv_1 _3789_ (.Y(_0377_),
    .A(net863));
 sg13g2_a22oi_1 _3790_ (.Y(_1727_),
    .B1(_1720_),
    .B2(net908),
    .A2(_0933_),
    .A1(net862));
 sg13g2_inv_1 _3791_ (.Y(_0378_),
    .A(net909));
 sg13g2_nor2b_1 _3792_ (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .B_N(_0056_),
    .Y(_1728_));
 sg13g2_o21ai_1 _3793_ (.B1(_0441_),
    .Y(_1729_),
    .A1(_0918_),
    .A2(_1728_));
 sg13g2_o21ai_1 _3794_ (.B1(_0936_),
    .Y(_1730_),
    .A1(_0441_),
    .A2(_0915_));
 sg13g2_nand2b_1 _3795_ (.Y(_1731_),
    .B(_1729_),
    .A_N(_1730_));
 sg13g2_o21ai_1 _3796_ (.B1(_1731_),
    .Y(_1732_),
    .A1(net360),
    .A2(_0942_));
 sg13g2_a22oi_1 _3797_ (.Y(_1733_),
    .B1(_1719_),
    .B2(_1732_),
    .A2(net579),
    .A1(net908));
 sg13g2_inv_1 _3798_ (.Y(_0379_),
    .A(_1733_));
 sg13g2_nand2_1 _3799_ (.Y(_1734_),
    .A(net360),
    .B(net579));
 sg13g2_o21ai_1 _3800_ (.B1(_0450_),
    .Y(_1735_),
    .A1(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .A2(net515));
 sg13g2_nand2_1 _3801_ (.Y(_1736_),
    .A(_0443_),
    .B(_0930_));
 sg13g2_o21ai_1 _3802_ (.B1(_1734_),
    .Y(_0380_),
    .A1(net516),
    .A2(_1736_));
 sg13g2_nor2_1 _3803_ (.A(_1961_),
    .B(_1980_),
    .Y(_1737_));
 sg13g2_nor3_2 _3804_ (.A(net342),
    .B(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ),
    .C(_1737_),
    .Y(_1738_));
 sg13g2_nor2_2 _3805_ (.A(net710),
    .B(_1738_),
    .Y(_1739_));
 sg13g2_nand2b_2 _3806_ (.Y(_1740_),
    .B(net740),
    .A_N(_1738_));
 sg13g2_nor2_1 _3807_ (.A(net318),
    .B(net600),
    .Y(_1741_));
 sg13g2_a21oi_1 _3808_ (.A1(net740),
    .A2(net318),
    .Y(_0381_),
    .B1(_1741_));
 sg13g2_a21oi_1 _3809_ (.A1(net318),
    .A2(net331),
    .Y(_1742_),
    .B1(_1738_));
 sg13g2_nor2_1 _3810_ (.A(net712),
    .B(_1742_),
    .Y(_1743_));
 sg13g2_a21oi_1 _3811_ (.A1(net740),
    .A2(net318),
    .Y(_1744_),
    .B1(net331));
 sg13g2_nor2_1 _3812_ (.A(_1743_),
    .B(_1744_),
    .Y(_0382_));
 sg13g2_o21ai_1 _3813_ (.B1(net202),
    .Y(_1745_),
    .A1(net712),
    .A2(_1742_));
 sg13g2_nand3_1 _3814_ (.B(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .C(net600),
    .A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .Y(_1746_));
 sg13g2_o21ai_1 _3815_ (.B1(_1745_),
    .Y(_0383_),
    .A1(net202),
    .A2(_1746_));
 sg13g2_and4_1 _3816_ (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .C(net202),
    .D(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .X(_1747_));
 sg13g2_o21ai_1 _3817_ (.B1(net740),
    .Y(_1748_),
    .A1(_1738_),
    .A2(_1747_));
 sg13g2_nand4_1 _3818_ (.B(net318),
    .C(net331),
    .A(net740),
    .Y(_1749_),
    .D(net202));
 sg13g2_nand2b_1 _3819_ (.Y(_1750_),
    .B(_1749_),
    .A_N(net1007));
 sg13g2_and2_1 _3820_ (.A(_1748_),
    .B(_1750_),
    .X(_0384_));
 sg13g2_nand2_1 _3821_ (.Y(_1751_),
    .A(net278),
    .B(_1748_));
 sg13g2_nand2_1 _3822_ (.Y(_1752_),
    .A(net600),
    .B(_1747_));
 sg13g2_o21ai_1 _3823_ (.B1(_1751_),
    .Y(_0385_),
    .A1(net278),
    .A2(_1752_));
 sg13g2_and3_2 _3824_ (.X(_1753_),
    .A(net278),
    .B(net287),
    .C(_1747_));
 sg13g2_nor2_1 _3825_ (.A(_1738_),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_nor2_1 _3826_ (.A(net712),
    .B(_1754_),
    .Y(_1755_));
 sg13g2_nand3_1 _3827_ (.B(net278),
    .C(_1747_),
    .A(net740),
    .Y(_1756_));
 sg13g2_a21oi_1 _3828_ (.A1(_1981_),
    .A2(_1756_),
    .Y(_0386_),
    .B1(_1755_));
 sg13g2_a21oi_1 _3829_ (.A1(net600),
    .A2(_1753_),
    .Y(_1757_),
    .B1(net172));
 sg13g2_a21oi_1 _3830_ (.A1(net172),
    .A2(_1755_),
    .Y(_0387_),
    .B1(_1757_));
 sg13g2_and3_1 _3831_ (.X(_1758_),
    .A(net172),
    .B(net873),
    .C(_1753_));
 sg13g2_a21oi_1 _3832_ (.A1(net172),
    .A2(_1753_),
    .Y(_1759_),
    .B1(net873));
 sg13g2_nor3_1 _3833_ (.A(_1740_),
    .B(_1758_),
    .C(_1759_),
    .Y(_1760_));
 sg13g2_a21o_1 _3834_ (.A2(net873),
    .A1(net710),
    .B1(_1760_),
    .X(_0388_));
 sg13g2_nand2_1 _3835_ (.Y(_1761_),
    .A(net710),
    .B(net402));
 sg13g2_and2_1 _3836_ (.A(net402),
    .B(_1758_),
    .X(_1762_));
 sg13g2_o21ai_1 _3837_ (.B1(net600),
    .Y(_1763_),
    .A1(net402),
    .A2(_1758_));
 sg13g2_o21ai_1 _3838_ (.B1(_1761_),
    .Y(_0389_),
    .A1(_1762_),
    .A2(_1763_));
 sg13g2_nand2_1 _3839_ (.Y(_1764_),
    .A(net710),
    .B(net393));
 sg13g2_and2_1 _3840_ (.A(net393),
    .B(_1762_),
    .X(_1765_));
 sg13g2_o21ai_1 _3841_ (.B1(_1739_),
    .Y(_1766_),
    .A1(net393),
    .A2(_1762_));
 sg13g2_o21ai_1 _3842_ (.B1(_1764_),
    .Y(_0390_),
    .A1(_1765_),
    .A2(_1766_));
 sg13g2_nand2_1 _3843_ (.Y(_1767_),
    .A(net710),
    .B(net303));
 sg13g2_and2_1 _3844_ (.A(net303),
    .B(_1765_),
    .X(_1768_));
 sg13g2_o21ai_1 _3845_ (.B1(net600),
    .Y(_1769_),
    .A1(net303),
    .A2(_1765_));
 sg13g2_o21ai_1 _3846_ (.B1(_1767_),
    .Y(_0391_),
    .A1(_1768_),
    .A2(_1769_));
 sg13g2_nand2_1 _3847_ (.Y(_1770_),
    .A(net710),
    .B(net422));
 sg13g2_xnor2_1 _3848_ (.Y(_1771_),
    .A(net422),
    .B(_1768_));
 sg13g2_o21ai_1 _3849_ (.B1(_1770_),
    .Y(_0392_),
    .A1(_1740_),
    .A2(_1771_));
 sg13g2_a21oi_1 _3850_ (.A1(net422),
    .A2(_1768_),
    .Y(_1772_),
    .B1(net887));
 sg13g2_and3_1 _3851_ (.X(_1773_),
    .A(net422),
    .B(net887),
    .C(_1768_));
 sg13g2_nor3_1 _3852_ (.A(_1740_),
    .B(_1772_),
    .C(_1773_),
    .Y(_1774_));
 sg13g2_a21o_1 _3853_ (.A2(net887),
    .A1(net710),
    .B1(_1774_),
    .X(_0393_));
 sg13g2_nand2_1 _3854_ (.Y(_1775_),
    .A(net710),
    .B(net366));
 sg13g2_and2_1 _3855_ (.A(net366),
    .B(_1773_),
    .X(_1776_));
 sg13g2_o21ai_1 _3856_ (.B1(net600),
    .Y(_1777_),
    .A1(net366),
    .A2(_1773_));
 sg13g2_o21ai_1 _3857_ (.B1(_1775_),
    .Y(_0394_),
    .A1(_1776_),
    .A2(_1777_));
 sg13g2_nand2_1 _3858_ (.Y(_1778_),
    .A(net711),
    .B(net297));
 sg13g2_and2_1 _3859_ (.A(net297),
    .B(_1776_),
    .X(_1779_));
 sg13g2_o21ai_1 _3860_ (.B1(_1739_),
    .Y(_1780_),
    .A1(net297),
    .A2(_1776_));
 sg13g2_o21ai_1 _3861_ (.B1(_1778_),
    .Y(_0395_),
    .A1(_1779_),
    .A2(_1780_));
 sg13g2_nand2_1 _3862_ (.Y(_1781_),
    .A(net711),
    .B(net305));
 sg13g2_and2_1 _3863_ (.A(net305),
    .B(_1779_),
    .X(_1782_));
 sg13g2_o21ai_1 _3864_ (.B1(_1739_),
    .Y(_1783_),
    .A1(net305),
    .A2(_1779_));
 sg13g2_o21ai_1 _3865_ (.B1(_1781_),
    .Y(_0396_),
    .A1(_1782_),
    .A2(_1783_));
 sg13g2_nand2_1 _3866_ (.Y(_1784_),
    .A(net711),
    .B(net566));
 sg13g2_nor2_1 _3867_ (.A(net566),
    .B(_1782_),
    .Y(_1785_));
 sg13g2_a21o_1 _3868_ (.A2(_1782_),
    .A1(net566),
    .B1(_1740_),
    .X(_1786_));
 sg13g2_a21oi_1 _3869_ (.A1(_1784_),
    .A2(_1786_),
    .Y(_0397_),
    .B1(_1785_));
 sg13g2_nand3_1 _3870_ (.B(net600),
    .C(_1782_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .Y(_1787_));
 sg13g2_a22oi_1 _3871_ (.Y(_0398_),
    .B1(_1787_),
    .B2(_1959_),
    .A2(_1786_),
    .A1(_0947_));
 sg13g2_a21oi_2 _3872_ (.B1(_0934_),
    .Y(_1788_),
    .A2(_0937_),
    .A1(_0935_));
 sg13g2_mux2_1 _3873_ (.A0(_1788_),
    .A1(net704),
    .S(net994),
    .X(_0399_));
 sg13g2_and2_1 _3874_ (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .B(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .X(_1789_));
 sg13g2_nand2_1 _3875_ (.Y(_1790_),
    .A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .B(net294));
 sg13g2_a21oi_1 _3876_ (.A1(_1788_),
    .A2(_1790_),
    .Y(_1791_),
    .B1(net704));
 sg13g2_a21oi_1 _3877_ (.A1(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .A2(_1788_),
    .Y(_1792_),
    .B1(net294));
 sg13g2_nor2_1 _3878_ (.A(_1791_),
    .B(net295),
    .Y(_0400_));
 sg13g2_a21oi_1 _3879_ (.A1(_1788_),
    .A2(_1789_),
    .Y(_1793_),
    .B1(net52));
 sg13g2_a21oi_1 _3880_ (.A1(net52),
    .A2(_1791_),
    .Y(_0401_),
    .B1(_1793_));
 sg13g2_nor2_1 _3881_ (.A(net712),
    .B(_1737_),
    .Y(_1794_));
 sg13g2_a21oi_1 _3882_ (.A1(net742),
    .A2(net287),
    .Y(_1795_),
    .B1(net878));
 sg13g2_nor2_1 _3883_ (.A(_1794_),
    .B(_1795_),
    .Y(_0402_));
 sg13g2_nor2_1 _3884_ (.A(net357),
    .B(net743),
    .Y(_1796_));
 sg13g2_a21oi_1 _3885_ (.A1(net741),
    .A2(_0975_),
    .Y(_0403_),
    .B1(net358));
 sg13g2_nor2_1 _3886_ (.A(net748),
    .B(net741),
    .Y(_1797_));
 sg13g2_a21oi_1 _3887_ (.A1(net741),
    .A2(net264),
    .Y(_0404_),
    .B1(_1797_));
 sg13g2_nor3_2 _3888_ (.A(_1961_),
    .B(net382),
    .C(net703),
    .Y(_1798_));
 sg13g2_o21ai_1 _3889_ (.B1(_1798_),
    .Y(_1799_),
    .A1(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .A2(net346));
 sg13g2_o21ai_1 _3890_ (.B1(_1799_),
    .Y(_0405_),
    .A1(_1937_),
    .A2(_0448_));
 sg13g2_nor2_1 _3891_ (.A(net746),
    .B(net743),
    .Y(_1800_));
 sg13g2_a21oi_1 _3892_ (.A1(net744),
    .A2(_0973_),
    .Y(_0406_),
    .B1(net977));
 sg13g2_mux2_1 _3893_ (.A0(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .A1(net973),
    .S(net704),
    .X(_0407_));
 sg13g2_nor2_1 _3894_ (.A(net913),
    .B(_0448_),
    .Y(_1801_));
 sg13g2_a21oi_1 _3895_ (.A1(_1935_),
    .A2(_0448_),
    .Y(_0408_),
    .B1(_1801_));
 sg13g2_mux2_1 _3896_ (.A0(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .A1(net852),
    .S(_0448_),
    .X(_0409_));
 sg13g2_nor2_1 _3897_ (.A(net386),
    .B(net703),
    .Y(_1802_));
 sg13g2_a21oi_1 _3898_ (.A1(_1935_),
    .A2(net704),
    .Y(_0410_),
    .B1(net387));
 sg13g2_o21ai_1 _3899_ (.B1(_1013_),
    .Y(_0411_),
    .A1(_1909_),
    .A2(net744));
 sg13g2_mux2_1 _3900_ (.A0(net967),
    .A1(net531),
    .S(net599),
    .X(_0412_));
 sg13g2_mux2_1 _3901_ (.A0(net940),
    .A1(net485),
    .S(net599),
    .X(_0413_));
 sg13g2_mux2_1 _3902_ (.A0(net945),
    .A1(net899),
    .S(net599),
    .X(_0414_));
 sg13g2_mux2_1 _3903_ (.A0(net966),
    .A1(net527),
    .S(net599),
    .X(_0415_));
 sg13g2_mux2_1 _3904_ (.A0(net929),
    .A1(net428),
    .S(_0972_),
    .X(_0416_));
 sg13g2_mux2_1 _3905_ (.A0(net992),
    .A1(net862),
    .S(_0972_),
    .X(_0417_));
 sg13g2_mux2_1 _3906_ (.A0(net982),
    .A1(net908),
    .S(net599),
    .X(_0418_));
 sg13g2_nor2_1 _3907_ (.A(\u_usb_cdc.u_sie.rx_data[7] ),
    .B(net599),
    .Y(_1803_));
 sg13g2_a21oi_1 _3908_ (.A1(net360),
    .A2(net599),
    .Y(_0419_),
    .B1(_1803_));
 sg13g2_nor2_1 _3909_ (.A(net735),
    .B(net234),
    .Y(_1804_));
 sg13g2_a21oi_1 _3910_ (.A1(net735),
    .A2(_0952_),
    .Y(_0420_),
    .B1(net235));
 sg13g2_nand2_1 _3911_ (.Y(_1805_),
    .A(net829),
    .B(_2003_));
 sg13g2_a22oi_1 _3912_ (.Y(_1806_),
    .B1(_0585_),
    .B2(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .A2(_2003_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ));
 sg13g2_nand2_1 _3913_ (.Y(_1807_),
    .A(_1805_),
    .B(_1806_));
 sg13g2_nor2_1 _3914_ (.A(net748),
    .B(net702),
    .Y(_1808_));
 sg13g2_a22oi_1 _3915_ (.Y(_1809_),
    .B1(_1952_),
    .B2(net831),
    .A2(_1938_),
    .A1(net838));
 sg13g2_a22oi_1 _3916_ (.Y(_1810_),
    .B1(\u_usb_cdc.u_sie.data_q[0] ),
    .B2(net835),
    .A2(\u_usb_cdc.u_sie.pid_q[0] ),
    .A1(net830));
 sg13g2_nand3_1 _3917_ (.B(_1809_),
    .C(_1810_),
    .A(_1696_),
    .Y(_1811_));
 sg13g2_a21o_1 _3918_ (.A2(_1811_),
    .A1(_1808_),
    .B1(_1807_),
    .X(_1812_));
 sg13g2_o21ai_1 _3919_ (.B1(_1812_),
    .Y(_1813_),
    .A1(net282),
    .A2(net705));
 sg13g2_nor2_1 _3920_ (.A(_1994_),
    .B(_1034_),
    .Y(_1814_));
 sg13g2_a21oi_1 _3921_ (.A1(net282),
    .A2(_1814_),
    .Y(_1815_),
    .B1(net622));
 sg13g2_a22oi_1 _3922_ (.Y(_0421_),
    .B1(_1813_),
    .B2(_1815_),
    .A2(net622),
    .A1(_1975_));
 sg13g2_nand2_1 _3923_ (.Y(_1816_),
    .A(net282),
    .B(net621));
 sg13g2_nor2_1 _3924_ (.A(_2003_),
    .B(net702),
    .Y(_1817_));
 sg13g2_nand2_2 _3925_ (.Y(_1818_),
    .A(net705),
    .B(_1034_));
 sg13g2_and2_1 _3926_ (.A(net705),
    .B(_1034_),
    .X(_1819_));
 sg13g2_a22oi_1 _3927_ (.Y(_1820_),
    .B1(_1939_),
    .B2(net838),
    .A2(\u_usb_cdc.u_sie.pid_q[1] ),
    .A1(net830));
 sg13g2_a22oi_1 _3928_ (.Y(_1821_),
    .B1(_1953_),
    .B2(net831),
    .A2(net765),
    .A1(net834));
 sg13g2_nand3_1 _3929_ (.B(_1820_),
    .C(_1821_),
    .A(_1991_),
    .Y(_1822_));
 sg13g2_a22oi_1 _3930_ (.Y(_1823_),
    .B1(_1822_),
    .B2(_1817_),
    .A2(_1818_),
    .A1(net211));
 sg13g2_a21oi_2 _3931_ (.B1(_1999_),
    .Y(_1824_),
    .A2(_1033_),
    .A1(net702));
 sg13g2_o21ai_1 _3932_ (.B1(net623),
    .Y(_1825_),
    .A1(_1993_),
    .A2(_1034_));
 sg13g2_nand2_1 _3933_ (.Y(_1826_),
    .A(_2005_),
    .B(_1824_));
 sg13g2_o21ai_1 _3934_ (.B1(_1816_),
    .Y(_0422_),
    .A1(_1823_),
    .A2(_1826_));
 sg13g2_nand2_1 _3935_ (.Y(_1827_),
    .A(net211),
    .B(net621));
 sg13g2_nand3_1 _3936_ (.B(\u_usb_cdc.ctrl_stall ),
    .C(_0572_),
    .A(net839),
    .Y(_1828_));
 sg13g2_a22oi_1 _3937_ (.Y(_1829_),
    .B1(net762),
    .B2(net834),
    .A2(\u_usb_cdc.u_sie.pid_q[2] ),
    .A1(net830));
 sg13g2_a22oi_1 _3938_ (.Y(_1830_),
    .B1(_1950_),
    .B2(net831),
    .A2(_1940_),
    .A1(net838));
 sg13g2_and3_1 _3939_ (.X(_1831_),
    .A(_1828_),
    .B(_1829_),
    .C(_1830_));
 sg13g2_o21ai_1 _3940_ (.B1(_1819_),
    .Y(_1832_),
    .A1(net702),
    .A2(_1831_));
 sg13g2_o21ai_1 _3941_ (.B1(_1832_),
    .Y(_1833_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.data_q[3] ),
    .A2(_1819_));
 sg13g2_o21ai_1 _3942_ (.B1(_1827_),
    .Y(_0423_),
    .A1(_1826_),
    .A2(_1833_));
 sg13g2_o21ai_1 _3943_ (.B1(_1990_),
    .Y(_1834_),
    .A1(_0579_),
    .A2(_1018_));
 sg13g2_a22oi_1 _3944_ (.Y(_1835_),
    .B1(_1951_),
    .B2(net831),
    .A2(_1941_),
    .A1(net838));
 sg13g2_a22oi_1 _3945_ (.Y(_1836_),
    .B1(\u_usb_cdc.u_sie.data_q[3] ),
    .B2(net834),
    .A2(\u_usb_cdc.u_sie.pid_q[3] ),
    .A1(net830));
 sg13g2_nand3_1 _3946_ (.B(_1835_),
    .C(_1836_),
    .A(_1834_),
    .Y(_1837_));
 sg13g2_nand2b_1 _3947_ (.Y(_1838_),
    .B(_2004_),
    .A_N(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ));
 sg13g2_o21ai_1 _3948_ (.B1(_1838_),
    .Y(_1839_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .A2(_2002_));
 sg13g2_nor2_1 _3949_ (.A(net702),
    .B(_1839_),
    .Y(_1840_));
 sg13g2_o21ai_1 _3950_ (.B1(_1840_),
    .Y(_1841_),
    .A1(_0585_),
    .A2(_1837_));
 sg13g2_o21ai_1 _3951_ (.B1(_1805_),
    .Y(_1842_),
    .A1(_1994_),
    .A2(_1034_));
 sg13g2_a21oi_1 _3952_ (.A1(\u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .A2(_1842_),
    .Y(_1843_),
    .B1(net621));
 sg13g2_a22oi_1 _3953_ (.Y(_0424_),
    .B1(_1841_),
    .B2(_1843_),
    .A2(net621),
    .A1(_1976_));
 sg13g2_nand2_1 _3954_ (.Y(_1844_),
    .A(_1990_),
    .B(_0579_));
 sg13g2_a22oi_1 _3955_ (.Y(_1845_),
    .B1(_1948_),
    .B2(net831),
    .A2(\u_usb_cdc.u_sie.data_q[4] ),
    .A1(net834));
 sg13g2_a22oi_1 _3956_ (.Y(_1846_),
    .B1(_1942_),
    .B2(\u_usb_cdc.u_sie.phy_state_q[4] ),
    .A2(_1922_),
    .A1(net830));
 sg13g2_nand3_1 _3957_ (.B(_1845_),
    .C(_1846_),
    .A(_1844_),
    .Y(_1847_));
 sg13g2_a21o_1 _3958_ (.A2(_1847_),
    .A1(_1808_),
    .B1(_1807_),
    .X(_1848_));
 sg13g2_o21ai_1 _3959_ (.B1(_1848_),
    .Y(_1849_),
    .A1(net274),
    .A2(net705));
 sg13g2_a21oi_1 _3960_ (.A1(net274),
    .A2(_1814_),
    .Y(_1850_),
    .B1(net622));
 sg13g2_a22oi_1 _3961_ (.Y(_0425_),
    .B1(_1849_),
    .B2(_1850_),
    .A2(net621),
    .A1(_1977_));
 sg13g2_nand2_1 _3962_ (.Y(_1851_),
    .A(net274),
    .B(net621));
 sg13g2_a22oi_1 _3963_ (.Y(_1852_),
    .B1(_1949_),
    .B2(net831),
    .A2(_1943_),
    .A1(net838));
 sg13g2_a22oi_1 _3964_ (.Y(_1853_),
    .B1(\u_usb_cdc.u_sie.data_q[5] ),
    .B2(net835),
    .A2(_1923_),
    .A1(net830));
 sg13g2_nand2_1 _3965_ (.Y(_1854_),
    .A(_1852_),
    .B(_1853_));
 sg13g2_a221oi_1 _3966_ (.B2(_1854_),
    .C1(_1818_),
    .B1(_1808_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .Y(_1855_),
    .A2(_0585_));
 sg13g2_o21ai_1 _3967_ (.B1(_1824_),
    .Y(_1856_),
    .A1(\u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .A2(_1819_));
 sg13g2_o21ai_1 _3968_ (.B1(_1851_),
    .Y(_0426_),
    .A1(_1855_),
    .A2(_1856_));
 sg13g2_a22oi_1 _3969_ (.Y(_1857_),
    .B1(_1947_),
    .B2(net831),
    .A2(_1924_),
    .A1(net830));
 sg13g2_a22oi_1 _3970_ (.Y(_1858_),
    .B1(\u_usb_cdc.u_sie.data_q[6] ),
    .B2(net834),
    .A2(_1944_),
    .A1(net838));
 sg13g2_nand3_1 _3971_ (.B(_1857_),
    .C(_1858_),
    .A(_0895_),
    .Y(_1859_));
 sg13g2_a21oi_1 _3972_ (.A1(_1808_),
    .A2(_1859_),
    .Y(_1860_),
    .B1(_1818_));
 sg13g2_a22oi_1 _3973_ (.Y(_1861_),
    .B1(_1860_),
    .B2(_1806_),
    .A2(_1818_),
    .A1(net368));
 sg13g2_a22oi_1 _3974_ (.Y(_1862_),
    .B1(_1824_),
    .B2(_1861_),
    .A2(net621),
    .A1(net400));
 sg13g2_inv_1 _3975_ (.Y(_0427_),
    .A(net401));
 sg13g2_or2_1 _3976_ (.X(_1863_),
    .B(_1696_),
    .A(_1018_));
 sg13g2_a22oi_1 _3977_ (.Y(_1864_),
    .B1(_1946_),
    .B2(net259),
    .A2(\u_usb_cdc.u_sie.data_q[7] ),
    .A1(net834));
 sg13g2_a22oi_1 _3978_ (.Y(_1865_),
    .B1(_1945_),
    .B2(\u_usb_cdc.u_sie.phy_state_q[4] ),
    .A2(_1925_),
    .A1(net830));
 sg13g2_nand4_1 _3979_ (.B(_1863_),
    .C(_1864_),
    .A(_1993_),
    .Y(_1866_),
    .D(_1865_));
 sg13g2_a221oi_1 _3980_ (.B2(_1866_),
    .C1(_1825_),
    .B1(_1817_),
    .A1(net829),
    .Y(_1867_),
    .A2(net705));
 sg13g2_a21o_1 _3981_ (.A2(net622),
    .A1(net368),
    .B1(_1867_),
    .X(_0428_));
 sg13g2_nor2_1 _3982_ (.A(net210),
    .B(_1824_),
    .Y(_1868_));
 sg13g2_a21oi_1 _3983_ (.A1(net210),
    .A2(net623),
    .Y(_0429_),
    .B1(_1868_));
 sg13g2_a21oi_1 _3984_ (.A1(net210),
    .A2(net623),
    .Y(_1869_),
    .B1(net312));
 sg13g2_o21ai_1 _3985_ (.B1(_2001_),
    .Y(_1870_),
    .A1(_1993_),
    .A2(_1034_));
 sg13g2_a21oi_1 _3986_ (.A1(_1998_),
    .A2(_1870_),
    .Y(_0430_),
    .B1(_1869_));
 sg13g2_xor2_1 _3987_ (.B(_2001_),
    .A(net1000),
    .X(_1871_));
 sg13g2_nor4_1 _3988_ (.A(net931),
    .B(_1999_),
    .C(_2003_),
    .D(_0954_),
    .Y(_1872_));
 sg13g2_a22oi_1 _3989_ (.Y(_1873_),
    .B1(_1033_),
    .B2(_1872_),
    .A2(net622),
    .A1(net1000));
 sg13g2_o21ai_1 _3990_ (.B1(net1001),
    .Y(_0431_),
    .A1(_1825_),
    .A2(_1871_));
 sg13g2_nand3_1 _3991_ (.B(_0440_),
    .C(_0917_),
    .A(net741),
    .Y(_1874_));
 sg13g2_o21ai_1 _3992_ (.B1(_1874_),
    .Y(_0432_),
    .A1(net741),
    .A2(_1980_));
 sg13g2_nand2b_1 _3993_ (.Y(_1875_),
    .B(_0586_),
    .A_N(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ));
 sg13g2_nand4_1 _3994_ (.B(net623),
    .C(_1838_),
    .A(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .Y(_1876_),
    .D(_1875_));
 sg13g2_nand2_1 _3995_ (.Y(_1877_),
    .A(net327),
    .B(net713));
 sg13g2_o21ai_1 _3996_ (.B1(_1877_),
    .Y(_0433_),
    .A1(net327),
    .A2(_1876_));
 sg13g2_nand2_1 _3997_ (.Y(_1878_),
    .A(net316),
    .B(net713));
 sg13g2_nand2_1 _3998_ (.Y(_1879_),
    .A(net327),
    .B(net316));
 sg13g2_xnor2_1 _3999_ (.Y(_1880_),
    .A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .B(net316));
 sg13g2_o21ai_1 _4000_ (.B1(_1878_),
    .Y(_0434_),
    .A1(_1876_),
    .A2(_1880_));
 sg13g2_nand2_1 _4001_ (.Y(_1881_),
    .A(net333),
    .B(net713));
 sg13g2_xor2_1 _4002_ (.B(_1879_),
    .A(net333),
    .X(_1882_));
 sg13g2_o21ai_1 _4003_ (.B1(_1881_),
    .Y(_0435_),
    .A1(_1876_),
    .A2(_1882_));
 sg13g2_o21ai_1 _4004_ (.B1(net624),
    .Y(_1883_),
    .A1(_1910_),
    .A2(_0612_));
 sg13g2_nor2_1 _4005_ (.A(net594),
    .B(_1883_),
    .Y(_1884_));
 sg13g2_nand2_1 _4006_ (.Y(_1885_),
    .A(net632),
    .B(_1884_));
 sg13g2_nand2_1 _4007_ (.Y(_1886_),
    .A(net85),
    .B(_1885_));
 sg13g2_o21ai_1 _4008_ (.B1(_1886_),
    .Y(_0436_),
    .A1(_1910_),
    .A2(_1885_));
 sg13g2_nand2_1 _4009_ (.Y(_1887_),
    .A(net634),
    .B(_1884_));
 sg13g2_nand2_1 _4010_ (.Y(_1888_),
    .A(net165),
    .B(_1887_));
 sg13g2_o21ai_1 _4011_ (.B1(_1888_),
    .Y(_0437_),
    .A1(_1910_),
    .A2(_1887_));
 sg13g2_mux2_1 _4012_ (.A0(_1041_),
    .A1(net828),
    .S(_1054_),
    .X(_1889_));
 sg13g2_mux2_1 _4013_ (.A0(net903),
    .A1(_1889_),
    .S(_1123_),
    .X(_0438_));
 sg13g2_nand2_1 _4014_ (.Y(_1890_),
    .A(net542),
    .B(_1054_));
 sg13g2_nand3_1 _4015_ (.B(net638),
    .C(_1890_),
    .A(net736),
    .Y(_1891_));
 sg13g2_o21ai_1 _4016_ (.B1(_1891_),
    .Y(_1892_),
    .A1(net737),
    .A2(net564));
 sg13g2_inv_1 _4017_ (.Y(_0439_),
    .A(net565));
 sg13g2_buf_1 _4018_ (.A(_0053_),
    .X(net37));
 sg13g2_dfrbpq_1 _4019_ (.RESET_B(net686),
    .D(net171),
    .Q(\u_usb_cdc.u_sie.out_toggle_q[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _4020_ (.RESET_B(net666),
    .D(net861),
    .Q(_0048_),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _4021_ (.RESET_B(net677),
    .D(net869),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _4022_ (.RESET_B(net666),
    .D(_0003_),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _4023_ (.RESET_B(net667),
    .D(net954),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _4024_ (.RESET_B(net676),
    .D(net972),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _4025_ (.RESET_B(net677),
    .D(_0006_),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _4026_ (.RESET_B(net676),
    .D(net907),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _4027_ (.RESET_B(net676),
    .D(net922),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _4028_ (.RESET_B(net666),
    .D(net846),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _4029_ (.RESET_B(net665),
    .D(net950),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _4030_ (.RESET_B(net665),
    .D(net207),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _4031_ (.RESET_B(net677),
    .D(net553),
    .Q(\u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _4032_ (.RESET_B(net689),
    .D(net851),
    .Q(\u_usb_cdc.u_sie.out_toggle_q[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _4033_ (.RESET_B(net691),
    .D(net311),
    .Q(\u_usb_cdc.u_sie.in_toggle_q[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _4034_ (.RESET_B(net681),
    .D(net925),
    .Q(\u_usb_cdc.u_sie.in_toggle_q[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _4035_ (.RESET_B(net681),
    .D(net356),
    .Q(\u_usb_cdc.u_sie.in_toggle_q[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _4036_ (.RESET_B(net678),
    .D(net537),
    .Q(_0049_),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4037_ (.RESET_B(net678),
    .D(net551),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _4038_ (.RESET_B(net678),
    .D(_0012_),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _4039_ (.RESET_B(net678),
    .D(net872),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4040_ (.RESET_B(net678),
    .D(net948),
    .Q(\u_usb_cdc.ctrl_stall ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _4041_ (.RESET_B(net678),
    .D(net867),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _4042_ (.RESET_B(net678),
    .D(net1004),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4043_ (.RESET_B(net685),
    .D(net889),
    .Q(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _4044_ (.RESET_B(net694),
    .D(net262),
    .Q(_0050_),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _4045_ (.RESET_B(net694),
    .D(net1051),
    .Q(\u_usb_cdc.u_sie.phy_state_q[1] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _4046_ (.RESET_B(net694),
    .D(net414),
    .Q(\u_usb_cdc.u_sie.phy_state_q[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _4047_ (.RESET_B(net694),
    .D(net526),
    .Q(\u_usb_cdc.u_sie.phy_state_q[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _4048_ (.RESET_B(net687),
    .D(_0023_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _4049_ (.RESET_B(net694),
    .D(net187),
    .Q(\u_usb_cdc.u_sie.phy_state_q[5] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _4050_ (.RESET_B(net697),
    .D(net209),
    .Q(\u_usb_cdc.u_sie.phy_state_q[6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _4051_ (.RESET_B(net687),
    .D(_0026_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[7] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4052_ (.RESET_B(net697),
    .D(net848),
    .Q(\u_usb_cdc.u_sie.phy_state_q[8] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _4053_ (.RESET_B(net694),
    .D(_0028_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _4054_ (.RESET_B(net695),
    .D(_0018_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4055_ (.RESET_B(net694),
    .D(_0019_),
    .Q(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _4056_ (.RESET_B(net731),
    .D(net353),
    .Q(_0051_),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _4057_ (.RESET_B(net728),
    .D(net893),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _4058_ (.RESET_B(net731),
    .D(net1013),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _4059_ (.RESET_B(net731),
    .D(_0031_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _4060_ (.RESET_B(net728),
    .D(net258),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _4061_ (.RESET_B(net724),
    .D(_0065_),
    .Q(_0052_),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _4062_ (.RESET_B(net724),
    .D(net344),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.state_q[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _4063_ (.RESET_B(net724),
    .D(_0034_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _4064_ (.RESET_B(net724),
    .D(_0035_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.state_q[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _4065_ (.RESET_B(net698),
    .D(net932),
    .Q(_0053_),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _4066_ (.RESET_B(net698),
    .D(net558),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _4067_ (.RESET_B(net698),
    .D(net383),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _4068_ (.RESET_B(net699),
    .D(_0038_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _4069_ (.RESET_B(net691),
    .D(net220),
    .Q(\u_usb_cdc.u_sie.addr_q[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _4070_ (.RESET_B(net699),
    .D(net309),
    .Q(_0054_),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _4071_ (.RESET_B(net672),
    .D(net543),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _4072_ (.RESET_B(net648),
    .D(_0075_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4073_ (.RESET_B(net652),
    .D(_0076_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4074_ (.RESET_B(net649),
    .D(_0077_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4075_ (.RESET_B(net648),
    .D(_0078_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4076_ (.RESET_B(net648),
    .D(_0079_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4077_ (.RESET_B(net650),
    .D(_0080_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4078_ (.RESET_B(net650),
    .D(_0081_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4079_ (.RESET_B(net650),
    .D(_0082_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _4080_ (.RESET_B(net654),
    .D(net379),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4081_ (.RESET_B(net649),
    .D(net443),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _4082_ (.RESET_B(net651),
    .D(net425),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4083_ (.RESET_B(net656),
    .D(net408),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4084_ (.RESET_B(net654),
    .D(net398),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4085_ (.RESET_B(net651),
    .D(net555),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4086_ (.RESET_B(net670),
    .D(net381),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4087_ (.RESET_B(net670),
    .D(net439),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4088_ (.RESET_B(net655),
    .D(net96),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4089_ (.RESET_B(net656),
    .D(net76),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4090_ (.RESET_B(net656),
    .D(net192),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4091_ (.RESET_B(net655),
    .D(net138),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4092_ (.RESET_B(net669),
    .D(net70),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4093_ (.RESET_B(net655),
    .D(net254),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4094_ (.RESET_B(net670),
    .D(net152),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4095_ (.RESET_B(net669),
    .D(net92),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4096_ (.RESET_B(net651),
    .D(net163),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4097_ (.RESET_B(net649),
    .D(net90),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4098_ (.RESET_B(net651),
    .D(net179),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4099_ (.RESET_B(net651),
    .D(net185),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4100_ (.RESET_B(net669),
    .D(net62),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4101_ (.RESET_B(net651),
    .D(net94),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4102_ (.RESET_B(net669),
    .D(net148),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4103_ (.RESET_B(net668),
    .D(net68),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _4104_ (.RESET_B(net649),
    .D(net419),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _4105_ (.RESET_B(net653),
    .D(net490),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _4106_ (.RESET_B(net656),
    .D(net427),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4107_ (.RESET_B(net656),
    .D(net453),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4108_ (.RESET_B(net671),
    .D(net482),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4109_ (.RESET_B(net656),
    .D(net411),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4110_ (.RESET_B(net669),
    .D(net457),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4111_ (.RESET_B(net668),
    .D(net474),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _4112_ (.RESET_B(net654),
    .D(net437),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4113_ (.RESET_B(net653),
    .D(net472),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4114_ (.RESET_B(net656),
    .D(net447),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4115_ (.RESET_B(net657),
    .D(net455),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4116_ (.RESET_B(net668),
    .D(net468),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4117_ (.RESET_B(net655),
    .D(net514),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4118_ (.RESET_B(net670),
    .D(net476),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4119_ (.RESET_B(net669),
    .D(net377),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4120_ (.RESET_B(net655),
    .D(net84),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4121_ (.RESET_B(net655),
    .D(net74),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4122_ (.RESET_B(net655),
    .D(net111),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4123_ (.RESET_B(net655),
    .D(net150),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _4124_ (.RESET_B(net669),
    .D(net131),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4125_ (.RESET_B(net657),
    .D(net57),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4126_ (.RESET_B(net670),
    .D(net72),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4127_ (.RESET_B(net669),
    .D(net81),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _4128_ (.RESET_B(net649),
    .D(net156),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4129_ (.RESET_B(net650),
    .D(net115),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4130_ (.RESET_B(net650),
    .D(net125),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4131_ (.RESET_B(net651),
    .D(net160),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4132_ (.RESET_B(net671),
    .D(net127),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4133_ (.RESET_B(net651),
    .D(net107),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4134_ (.RESET_B(net670),
    .D(net88),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _4135_ (.RESET_B(net670),
    .D(net60),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _4136_ (.RESET_B(net649),
    .D(net396),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _4137_ (.RESET_B(net648),
    .D(net435),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _4138_ (.RESET_B(net650),
    .D(net512),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4139_ (.RESET_B(net650),
    .D(net494),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4140_ (.RESET_B(net668),
    .D(net488),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _4141_ (.RESET_B(net650),
    .D(net484),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _4142_ (.RESET_B(net672),
    .D(net463),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _4143_ (.RESET_B(net668),
    .D(net338),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[63] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _4144_ (.RESET_B(net653),
    .D(net451),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4145_ (.RESET_B(net653),
    .D(net431),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _4146_ (.RESET_B(net653),
    .D(net465),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _4147_ (.RESET_B(net654),
    .D(net478),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _4148_ (.RESET_B(net668),
    .D(net449),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4149_ (.RESET_B(net654),
    .D(net433),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4150_ (.RESET_B(net674),
    .D(net470),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _4151_ (.RESET_B(net674),
    .D(net492),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[71] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _4152_ (.RESET_B(net683),
    .D(_0155_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _4153_ (.RESET_B(net683),
    .D(_0156_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _4154_ (.RESET_B(net683),
    .D(net902),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _4155_ (.RESET_B(net648),
    .D(_0158_),
    .Q(\u_usb_cdc.in_ready_o [0]),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _4156_ (.RESET_B(net672),
    .D(net998),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4157_ (.RESET_B(net672),
    .D(_0160_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _4158_ (.RESET_B(net672),
    .D(_0161_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4159_ (.RESET_B(net672),
    .D(_0162_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _4160_ (.RESET_B(net673),
    .D(net302),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4161_ (.RESET_B(net672),
    .D(net928),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _4162_ (.RESET_B(net673),
    .D(net281),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4163_ (.RESET_B(net673),
    .D(net336),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _4164_ (.RESET_B(net665),
    .D(net256),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4165_ (.RESET_B(net661),
    .D(_0168_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _4166_ (.RESET_B(net659),
    .D(_0169_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4167_ (.RESET_B(net644),
    .D(_0170_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4168_ (.RESET_B(net661),
    .D(net158),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4169_ (.RESET_B(net663),
    .D(net233),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4170_ (.RESET_B(net644),
    .D(net55),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4171_ (.RESET_B(net662),
    .D(_0174_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4172_ (.RESET_B(net660),
    .D(net105),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4173_ (.RESET_B(net660),
    .D(net217),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4174_ (.RESET_B(net645),
    .D(net123),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4175_ (.RESET_B(net644),
    .D(net103),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[11] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4176_ (.RESET_B(net659),
    .D(net154),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4177_ (.RESET_B(net662),
    .D(net226),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4178_ (.RESET_B(net647),
    .D(net181),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[14] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4179_ (.RESET_B(net646),
    .D(net222),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4180_ (.RESET_B(net645),
    .D(net390),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4181_ (.RESET_B(net645),
    .D(net547),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _4182_ (.RESET_B(net645),
    .D(net322),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[18] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4183_ (.RESET_B(net639),
    .D(net441),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _4184_ (.RESET_B(net647),
    .D(net300),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4185_ (.RESET_B(net646),
    .D(net284),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4186_ (.RESET_B(net645),
    .D(net268),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4187_ (.RESET_B(net646),
    .D(net315),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[23] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4188_ (.RESET_B(net665),
    .D(net228),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4189_ (.RESET_B(net665),
    .D(_0192_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _4190_ (.RESET_B(net661),
    .D(_0193_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[26] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4191_ (.RESET_B(net644),
    .D(_0194_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4192_ (.RESET_B(net661),
    .D(net177),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[28] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _4193_ (.RESET_B(net663),
    .D(net205),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[29] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _4194_ (.RESET_B(net645),
    .D(net183),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4195_ (.RESET_B(net662),
    .D(_0198_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[31] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4196_ (.RESET_B(net665),
    .D(net243),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _4197_ (.RESET_B(net661),
    .D(_0200_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _4198_ (.RESET_B(net659),
    .D(_0201_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4199_ (.RESET_B(net644),
    .D(_0202_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[35] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4200_ (.RESET_B(net664),
    .D(net241),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4201_ (.RESET_B(net662),
    .D(net99),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4202_ (.RESET_B(net644),
    .D(net140),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[38] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4203_ (.RESET_B(net662),
    .D(net142),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4204_ (.RESET_B(net659),
    .D(net79),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4205_ (.RESET_B(net659),
    .D(net247),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4206_ (.RESET_B(net645),
    .D(net133),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _4207_ (.RESET_B(net644),
    .D(net196),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4208_ (.RESET_B(net660),
    .D(net65),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4209_ (.RESET_B(net662),
    .D(net109),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4210_ (.RESET_B(net646),
    .D(net198),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4211_ (.RESET_B(net647),
    .D(net113),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4212_ (.RESET_B(net659),
    .D(net363),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4213_ (.RESET_B(net659),
    .D(net417),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4214_ (.RESET_B(net647),
    .D(net277),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4215_ (.RESET_B(net639),
    .D(net326),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[51] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _4216_ (.RESET_B(net660),
    .D(net324),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _4217_ (.RESET_B(net642),
    .D(net501),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4218_ (.RESET_B(net642),
    .D(net330),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[54] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _4219_ (.RESET_B(net646),
    .D(net273),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _4220_ (.RESET_B(net665),
    .D(net224),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _4221_ (.RESET_B(net661),
    .D(_0224_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _4222_ (.RESET_B(net659),
    .D(_0225_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4223_ (.RESET_B(net644),
    .D(_0226_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[59] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _4224_ (.RESET_B(net664),
    .D(net249),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _4225_ (.RESET_B(net663),
    .D(net168),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4226_ (.RESET_B(net646),
    .D(net129),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[62] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4227_ (.RESET_B(net662),
    .D(_0230_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4228_ (.RESET_B(net639),
    .D(net119),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[64] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4229_ (.RESET_B(net639),
    .D(net146),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[65] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _4230_ (.RESET_B(net639),
    .D(net121),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[66] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4231_ (.RESET_B(net639),
    .D(net194),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[67] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _4232_ (.RESET_B(net639),
    .D(net101),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[68] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4233_ (.RESET_B(net641),
    .D(net135),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[69] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4234_ (.RESET_B(net639),
    .D(net117),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[70] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4235_ (.RESET_B(net643),
    .D(net144),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[71] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4236_ (.RESET_B(net653),
    .D(_0239_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4237_ (.RESET_B(net646),
    .D(_0240_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _4238_ (.RESET_B(net646),
    .D(net1058),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _4239_ (.RESET_B(net642),
    .D(_0242_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4240_ (.RESET_B(net640),
    .D(net406),
    .Q(net29),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4241_ (.RESET_B(net640),
    .D(net895),
    .Q(net30),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _4242_ (.RESET_B(net640),
    .D(net496),
    .Q(net31),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4243_ (.RESET_B(net640),
    .D(net560),
    .Q(net32),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4244_ (.RESET_B(net640),
    .D(net545),
    .Q(net33),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _4245_ (.RESET_B(net640),
    .D(net898),
    .Q(net34),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _4246_ (.RESET_B(net640),
    .D(net877),
    .Q(net35),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _4247_ (.RESET_B(net640),
    .D(net875),
    .Q(net36),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4248_ (.RESET_B(net653),
    .D(net956),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4249_ (.RESET_B(net653),
    .D(net969),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4250_ (.RESET_B(net654),
    .D(net984),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4251_ (.RESET_B(net649),
    .D(net961),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _4252_ (.RESET_B(net641),
    .D(net534),
    .Q(\u_usb_cdc.out_valid_o [0]),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4253_ (.RESET_B(net643),
    .D(net1055),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _4254_ (.RESET_B(net642),
    .D(_0256_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _4255_ (.RESET_B(net642),
    .D(net1025),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _4256_ (.RESET_B(net643),
    .D(_0258_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _4257_ (.RESET_B(net683),
    .D(net1047),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _4258_ (.RESET_B(net683),
    .D(net1028),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4259_ (.RESET_B(net683),
    .D(net990),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _4260_ (.RESET_B(net673),
    .D(_0262_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _4261_ (.RESET_B(net676),
    .D(_0263_),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _4262_ (.RESET_B(net676),
    .D(_0264_),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _4263_ (.RESET_B(net676),
    .D(_0265_),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _4264_ (.RESET_B(net676),
    .D(_0266_),
    .Q(\u_usb_cdc.u_ctrl_endp.endp_q[3] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _4265_ (.RESET_B(net676),
    .D(net480),
    .Q(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _4266_ (.RESET_B(net679),
    .D(net270),
    .Q(\u_usb_cdc.addr[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _4267_ (.RESET_B(net680),
    .D(_0269_),
    .Q(\u_usb_cdc.addr[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _4268_ (.RESET_B(net693),
    .D(_0270_),
    .Q(\u_usb_cdc.addr[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _4269_ (.RESET_B(net679),
    .D(_0271_),
    .Q(\u_usb_cdc.addr[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _4270_ (.RESET_B(net693),
    .D(_0272_),
    .Q(\u_usb_cdc.addr[4] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _4271_ (.RESET_B(net693),
    .D(_0273_),
    .Q(\u_usb_cdc.addr[5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _4272_ (.RESET_B(net680),
    .D(_0274_),
    .Q(\u_usb_cdc.addr[6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _4273_ (.RESET_B(net679),
    .D(_0275_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _4274_ (.RESET_B(net679),
    .D(_0276_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _4275_ (.RESET_B(net693),
    .D(_0277_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _4276_ (.RESET_B(net679),
    .D(_0278_),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[3] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _4277_ (.RESET_B(net693),
    .D(net385),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[4] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _4278_ (.RESET_B(net693),
    .D(net459),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[5] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _4279_ (.RESET_B(net680),
    .D(net365),
    .Q(\u_usb_cdc.u_ctrl_endp.addr_dd[6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _4280_ (.RESET_B(net677),
    .D(_0282_),
    .Q(_0055_),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _4281_ (.RESET_B(net679),
    .D(_0283_),
    .Q(\u_usb_cdc.u_ctrl_endp.dev_state_q[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _4282_ (.RESET_B(net665),
    .D(_0284_),
    .Q(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _4283_ (.RESET_B(net677),
    .D(_0285_),
    .Q(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _4284_ (.RESET_B(net666),
    .D(net885),
    .Q(\u_usb_cdc.u_ctrl_endp.class_q ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _4285_ (.RESET_B(net677),
    .D(_0287_),
    .Q(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _4286_ (.RESET_B(net666),
    .D(_0288_),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4287_ (.RESET_B(net666),
    .D(_0289_),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4288_ (.RESET_B(net666),
    .D(net524),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4289_ (.RESET_B(net662),
    .D(net917),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _4290_ (.RESET_B(net663),
    .D(net539),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4291_ (.RESET_B(net663),
    .D(net855),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _4292_ (.RESET_B(net667),
    .D(net891),
    .Q(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4293_ (.RESET_B(net674),
    .D(_0295_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4294_ (.RESET_B(net674),
    .D(_0296_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _4295_ (.RESET_B(net674),
    .D(_0297_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4296_ (.RESET_B(net674),
    .D(_0298_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _4297_ (.RESET_B(net674),
    .D(_0299_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _4298_ (.RESET_B(net674),
    .D(_0300_),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _4299_ (.RESET_B(net668),
    .D(net952),
    .Q(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _4300_ (.RESET_B(net668),
    .D(_0302_),
    .Q(\u_usb_cdc.bulk_out_nak [0]),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _4301_ (.RESET_B(net686),
    .D(net943),
    .Q(\u_usb_cdc.endp[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _4302_ (.RESET_B(net681),
    .D(net959),
    .Q(\u_usb_cdc.endp[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _4303_ (.RESET_B(net691),
    .D(_0305_),
    .Q(\u_usb_cdc.endp[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _4304_ (.RESET_B(net691),
    .D(net965),
    .Q(\u_usb_cdc.endp[3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _4305_ (.RESET_B(net679),
    .D(_0307_),
    .Q(\u_usb_cdc.u_sie.addr_q[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _4306_ (.RESET_B(net693),
    .D(_0308_),
    .Q(\u_usb_cdc.u_sie.addr_q[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _4307_ (.RESET_B(net679),
    .D(_0309_),
    .Q(\u_usb_cdc.u_sie.addr_q[3] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _4308_ (.RESET_B(net691),
    .D(net238),
    .Q(\u_usb_cdc.u_sie.addr_q[4] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _4309_ (.RESET_B(net693),
    .D(net215),
    .Q(\u_usb_cdc.u_sie.addr_q[5] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _4310_ (.RESET_B(net680),
    .D(net251),
    .Q(\u_usb_cdc.u_sie.addr_q[6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _4311_ (.RESET_B(net734),
    .D(net938),
    .Q(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _4312_ (.RESET_B(net734),
    .D(net348),
    .Q(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _4313_ (.RESET_B(net686),
    .D(_0315_),
    .Q(\u_usb_cdc.sie_in_req ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4314_ (.RESET_B(net691),
    .D(net1006),
    .Q(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _4315_ (.RESET_B(net692),
    .D(net509),
    .Q(\u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _4316_ (.RESET_B(net692),
    .D(net461),
    .Q(\u_usb_cdc.u_sie.delay_cnt_q[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _4317_ (.RESET_B(net684),
    .D(net290),
    .Q(\u_usb_cdc.u_sie.in_byte_q[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _4318_ (.RESET_B(net683),
    .D(net320),
    .Q(\u_usb_cdc.u_sie.in_byte_q[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _4319_ (.RESET_B(net684),
    .D(net231),
    .Q(\u_usb_cdc.u_sie.in_byte_q[2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _4320_ (.RESET_B(net684),
    .D(net340),
    .Q(\u_usb_cdc.u_sie.in_byte_q[3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _4321_ (.RESET_B(net695),
    .D(_0323_),
    .Q(\u_usb_cdc.u_sie.crc16_q[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _4322_ (.RESET_B(net695),
    .D(_0324_),
    .Q(\u_usb_cdc.u_sie.crc16_q[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _4323_ (.RESET_B(net688),
    .D(_0325_),
    .Q(\u_usb_cdc.u_sie.crc16_q[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4324_ (.RESET_B(net688),
    .D(_0326_),
    .Q(\u_usb_cdc.u_sie.crc16_q[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4325_ (.RESET_B(net687),
    .D(_0327_),
    .Q(\u_usb_cdc.u_sie.crc16_q[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4326_ (.RESET_B(net687),
    .D(_0328_),
    .Q(\u_usb_cdc.u_sie.crc16_q[5] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4327_ (.RESET_B(net688),
    .D(_0329_),
    .Q(\u_usb_cdc.u_sie.crc16_q[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4328_ (.RESET_B(net688),
    .D(net883),
    .Q(\u_usb_cdc.u_sie.crc16_q[7] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4329_ (.RESET_B(net695),
    .D(_0331_),
    .Q(\u_usb_cdc.u_sie.crc16_q[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _4330_ (.RESET_B(net687),
    .D(_0332_),
    .Q(\u_usb_cdc.u_sie.crc16_q[9] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _4331_ (.RESET_B(net688),
    .D(_0333_),
    .Q(\u_usb_cdc.u_sie.crc16_q[10] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4332_ (.RESET_B(net687),
    .D(net373),
    .Q(\u_usb_cdc.u_sie.crc16_q[11] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _4333_ (.RESET_B(net687),
    .D(net286),
    .Q(\u_usb_cdc.u_sie.crc16_q[12] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _4334_ (.RESET_B(net687),
    .D(net307),
    .Q(\u_usb_cdc.u_sie.crc16_q[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _4335_ (.RESET_B(net695),
    .D(net350),
    .Q(\u_usb_cdc.u_sie.crc16_q[14] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _4336_ (.RESET_B(net695),
    .D(_0338_),
    .Q(\u_usb_cdc.u_sie.crc16_q[15] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4337_ (.RESET_B(net685),
    .D(_0339_),
    .Q(\u_usb_cdc.u_sie.data_q[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4338_ (.RESET_B(net685),
    .D(_0340_),
    .Q(\u_usb_cdc.u_sie.data_q[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _4339_ (.RESET_B(net685),
    .D(_0341_),
    .Q(\u_usb_cdc.u_sie.data_q[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _4340_ (.RESET_B(net686),
    .D(_0342_),
    .Q(\u_usb_cdc.u_sie.data_q[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4341_ (.RESET_B(net686),
    .D(_0343_),
    .Q(\u_usb_cdc.u_sie.data_q[4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4342_ (.RESET_B(net686),
    .D(_0344_),
    .Q(\u_usb_cdc.u_sie.data_q[5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4343_ (.RESET_B(net686),
    .D(_0345_),
    .Q(\u_usb_cdc.u_sie.data_q[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4344_ (.RESET_B(net686),
    .D(_0346_),
    .Q(\u_usb_cdc.u_sie.data_q[7] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4345_ (.RESET_B(net681),
    .D(_0347_),
    .Q(\u_usb_cdc.sie_out_data[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _4346_ (.RESET_B(net682),
    .D(_0348_),
    .Q(\u_usb_cdc.sie_out_data[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _4347_ (.RESET_B(net691),
    .D(_0349_),
    .Q(\u_usb_cdc.sie_out_data[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _4348_ (.RESET_B(net681),
    .D(_0350_),
    .Q(\u_usb_cdc.sie_out_data[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _4349_ (.RESET_B(net681),
    .D(_0351_),
    .Q(\u_usb_cdc.sie_out_data[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _4350_ (.RESET_B(net691),
    .D(_0352_),
    .Q(\u_usb_cdc.sie_out_data[5] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _4351_ (.RESET_B(net681),
    .D(_0353_),
    .Q(\u_usb_cdc.sie_out_data[6] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _4352_ (.RESET_B(net681),
    .D(_0354_),
    .Q(\u_usb_cdc.sie_out_data[7] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _4353_ (.RESET_B(net641),
    .D(_0355_),
    .Q(net14),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4354_ (.RESET_B(net641),
    .D(net421),
    .Q(net15),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _4355_ (.RESET_B(net641),
    .D(net375),
    .Q(net16),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4356_ (.RESET_B(net642),
    .D(net506),
    .Q(net17),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4357_ (.RESET_B(net642),
    .D(net859),
    .Q(net18),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _4358_ (.RESET_B(net648),
    .D(net371),
    .Q(net19),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _4359_ (.RESET_B(net648),
    .D(net504),
    .Q(net20),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _4360_ (.RESET_B(net648),
    .D(net844),
    .Q(net21),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _4361_ (.RESET_B(net641),
    .D(net912),
    .Q(net26),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4362_ (.RESET_B(net641),
    .D(net963),
    .Q(net27),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _4363_ (.RESET_B(net641),
    .D(net934),
    .Q(net28),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _4364_ (.RESET_B(net695),
    .D(_0366_),
    .Q(\u_usb_cdc.u_sie.pid_q[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4365_ (.RESET_B(net695),
    .D(_0367_),
    .Q(\u_usb_cdc.u_sie.pid_q[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4366_ (.RESET_B(net694),
    .D(net1010),
    .Q(\u_usb_cdc.u_sie.pid_q[2] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _4367_ (.RESET_B(net689),
    .D(net1019),
    .Q(\u_usb_cdc.u_sie.pid_q[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _4368_ (.RESET_B(net692),
    .D(_0370_),
    .Q(\u_usb_cdc.sie_out_err ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _4369_ (.RESET_B(net692),
    .D(net293),
    .Q(\u_usb_cdc.u_sie.out_eop_q ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _4370_ (.RESET_B(net728),
    .D(_0372_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _4371_ (.RESET_B(net728),
    .D(_0373_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _4372_ (.RESET_B(net729),
    .D(_0374_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _4373_ (.RESET_B(net730),
    .D(_0375_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _4374_ (.RESET_B(net730),
    .D(_0376_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _4375_ (.RESET_B(net730),
    .D(_0377_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _4376_ (.RESET_B(net730),
    .D(_0378_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _4377_ (.RESET_B(net730),
    .D(_0379_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _4378_ (.RESET_B(net732),
    .D(net517),
    .Q(_0056_),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _4379_ (.RESET_B(net723),
    .D(_0381_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _4380_ (.RESET_B(net722),
    .D(net332),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _4381_ (.RESET_B(net722),
    .D(net203),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _4382_ (.RESET_B(net722),
    .D(net1008),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _4383_ (.RESET_B(net722),
    .D(net279),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _4384_ (.RESET_B(net722),
    .D(net288),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _4385_ (.RESET_B(net722),
    .D(net173),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _4386_ (.RESET_B(net723),
    .D(_0388_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _4387_ (.RESET_B(net723),
    .D(net403),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _4388_ (.RESET_B(net723),
    .D(net394),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _4389_ (.RESET_B(net723),
    .D(net304),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _4390_ (.RESET_B(net722),
    .D(_0392_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _4391_ (.RESET_B(net726),
    .D(_0393_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _4392_ (.RESET_B(net726),
    .D(net367),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _4393_ (.RESET_B(net726),
    .D(net298),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _4394_ (.RESET_B(net726),
    .D(_0396_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _4395_ (.RESET_B(net726),
    .D(_0397_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _4396_ (.RESET_B(net725),
    .D(net190),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _4397_ (.RESET_B(net727),
    .D(_0399_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _4398_ (.RESET_B(net725),
    .D(net296),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _4399_ (.RESET_B(net725),
    .D(net53),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _4400_ (.RESET_B(net724),
    .D(net879),
    .Q(\u_usb_cdc.bus_reset ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _4401_ (.RESET_B(net728),
    .D(net359),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _4402_ (.RESET_B(net728),
    .D(_0404_),
    .Q(\u_usb_cdc.u_sie.rx_err ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _4403_ (.RESET_B(net725),
    .D(net936),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _4404_ (.RESET_B(net728),
    .D(_0043_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_q ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _4405_ (.RESET_B(net729),
    .D(net978),
    .Q(\u_usb_cdc.u_sie.rx_valid ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _4406_ (.RESET_B(net728),
    .D(_0044_),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_err_q ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _4407_ (.RESET_B(net731),
    .D(net974),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _4408_ (.RESET_B(net731),
    .D(net914),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _4409_ (.RESET_B(net727),
    .D(net853),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _4410_ (.RESET_B(net731),
    .D(net388),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _4411_ (.RESET_B(net685),
    .D(net1035),
    .Q(\u_usb_cdc.sie_in_data_ack ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _4412_ (.RESET_B(net729),
    .D(net530),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.rx_valid_q ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _4413_ (.RESET_B(net729),
    .D(_0412_),
    .Q(\u_usb_cdc.u_sie.rx_data[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _4414_ (.RESET_B(net729),
    .D(_0413_),
    .Q(\u_usb_cdc.u_sie.rx_data[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _4415_ (.RESET_B(net729),
    .D(_0414_),
    .Q(\u_usb_cdc.u_sie.rx_data[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _4416_ (.RESET_B(net729),
    .D(_0415_),
    .Q(\u_usb_cdc.u_sie.rx_data[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _4417_ (.RESET_B(net730),
    .D(net930),
    .Q(\u_usb_cdc.u_sie.rx_data[4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _4418_ (.RESET_B(net730),
    .D(_0417_),
    .Q(\u_usb_cdc.u_sie.rx_data[5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _4419_ (.RESET_B(net730),
    .D(_0418_),
    .Q(\u_usb_cdc.u_sie.rx_data[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _4420_ (.RESET_B(net729),
    .D(net361),
    .Q(\u_usb_cdc.u_sie.rx_data[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _4421_ (.RESET_B(net725),
    .D(net50),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _4422_ (.RESET_B(net725),
    .D(net522),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _4423_ (.RESET_B(net734),
    .D(net236),
    .Q(\u_usb_cdc.dp_pu_o ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _4424_ (.RESET_B(net727),
    .D(net47),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _4425_ (.RESET_B(net725),
    .D(net44),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _4426_ (.RESET_B(net725),
    .D(net13),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _4427_ (.RESET_B(net731),
    .D(net46),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _4428_ (.RESET_B(net732),
    .D(net43),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _4429_ (.RESET_B(net732),
    .D(net12),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _4430_ (.RESET_B(net699),
    .D(_0421_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _4431_ (.RESET_B(net698),
    .D(_0422_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _4432_ (.RESET_B(net696),
    .D(net212),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _4433_ (.RESET_B(net696),
    .D(net266),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _4434_ (.RESET_B(net698),
    .D(_0425_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _4435_ (.RESET_B(net696),
    .D(net275),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _4436_ (.RESET_B(net696),
    .D(_0427_),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _4437_ (.RESET_B(net696),
    .D(net369),
    .Q(_0057_),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _4438_ (.RESET_B(net698),
    .D(_0429_),
    .Q(_0058_),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _4439_ (.RESET_B(net698),
    .D(net313),
    .Q(_0059_),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _4440_ (.RESET_B(net698),
    .D(_0431_),
    .Q(_0060_),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _4441_ (.RESET_B(net724),
    .D(net245),
    .Q(\u_usb_cdc.u_sie.u_phy_rx.se0_q ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _4442_ (.RESET_B(net699),
    .D(net328),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _4443_ (.RESET_B(net699),
    .D(net317),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _4444_ (.RESET_B(net699),
    .D(net334),
    .Q(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _4445_ (.RESET_B(net726),
    .D(_0041_),
    .Q(\u_usb_cdc.clk_gate_q ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _4446_ (.RESET_B(net726),
    .D(_0039_),
    .Q(\u_usb_cdc.clk_cnt_q[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _4447_ (.RESET_B(net726),
    .D(_0040_),
    .Q(\u_usb_cdc.clk_cnt_q[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _4448_ (.RESET_B(net1),
    .D(net45),
    .Q(\u_usb_cdc.rstn ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4449_ (.RESET_B(net1),
    .D(net42),
    .Q(\u_usb_cdc.rstn_sq[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _4450_ (.RESET_B(net684),
    .D(net86),
    .Q(\u_usb_cdc.u_sie.in_zlp_q[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _4451_ (.RESET_B(net684),
    .D(net166),
    .Q(\u_usb_cdc.u_sie.in_zlp_q[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _4452_ (.RESET_B(net683),
    .D(_0438_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _4453_ (.RESET_B(net672),
    .D(_0439_),
    .Q(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _4449__42 (.L_HI(net42));
 sg13g2_buf_1 _4456_ (.A(\u_usb_cdc.out_valid_o [0]),
    .X(net22));
 sg13g2_buf_1 _4457_ (.A(\u_usb_cdc.in_ready_o [0]),
    .X(net23));
 sg13g2_buf_1 _4458_ (.A(\u_usb_cdc.dp_pu_o ),
    .X(net24));
 sg13g2_buf_8 _4459_ (.A(\u_usb_cdc.configured_o ),
    .X(net25));
 sg13g2_buf_1 _4460_ (.A(net37),
    .X(net39));
 sg13g2_buf_8 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_8 fanout568 (.A(_1406_),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(_1377_),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(_1388_),
    .X(net570));
 sg13g2_buf_1 fanout571 (.A(_1388_),
    .X(net571));
 sg13g2_buf_8 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_8 fanout573 (.A(_1484_),
    .X(net573));
 sg13g2_buf_8 fanout574 (.A(_0693_),
    .X(net574));
 sg13g2_buf_8 fanout575 (.A(net577),
    .X(net575));
 sg13g2_buf_1 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_8 fanout577 (.A(_1483_),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(_1254_),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(_0933_),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(net582),
    .X(net580));
 sg13g2_buf_1 fanout581 (.A(net582),
    .X(net581));
 sg13g2_buf_8 fanout582 (.A(_0869_),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(_0637_),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_0636_),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_1 fanout588 (.A(_0627_),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(_0602_),
    .X(net589));
 sg13g2_buf_8 fanout590 (.A(net592),
    .X(net590));
 sg13g2_buf_1 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(_0594_),
    .X(net592));
 sg13g2_buf_8 fanout593 (.A(net596),
    .X(net593));
 sg13g2_buf_8 fanout594 (.A(net596),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(net596),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(_0593_),
    .X(net596));
 sg13g2_buf_8 fanout597 (.A(_0592_),
    .X(net597));
 sg13g2_buf_8 fanout598 (.A(_0592_),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(_0972_),
    .X(net599));
 sg13g2_buf_8 fanout600 (.A(_1739_),
    .X(net600));
 sg13g2_buf_8 fanout601 (.A(_1275_),
    .X(net601));
 sg13g2_buf_1 fanout602 (.A(_1275_),
    .X(net602));
 sg13g2_buf_8 fanout603 (.A(_1119_),
    .X(net603));
 sg13g2_buf_8 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_8 fanout605 (.A(_1211_),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(_1193_),
    .X(net607));
 sg13g2_buf_8 fanout608 (.A(net610),
    .X(net608));
 sg13g2_buf_1 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(_1184_),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(_1166_),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(_1166_),
    .X(net612));
 sg13g2_buf_8 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(_1137_),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(_1099_),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(_1064_),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(_0711_),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(_0658_),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(_1999_),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(_1998_),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_1488_),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(_1360_),
    .X(net626));
 sg13g2_buf_8 fanout627 (.A(net629),
    .X(net627));
 sg13g2_buf_1 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(_1220_),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(_1135_),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_1 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(_0575_),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(_0572_),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(_0450_),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(_1061_),
    .X(net636));
 sg13g2_buf_8 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(_1038_),
    .X(net638));
 sg13g2_buf_8 fanout639 (.A(net643),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net643),
    .X(net640));
 sg13g2_buf_8 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_8 fanout643 (.A(net658),
    .X(net643));
 sg13g2_buf_8 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_8 fanout645 (.A(net647),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(net647),
    .X(net646));
 sg13g2_buf_8 fanout647 (.A(net658),
    .X(net647));
 sg13g2_buf_8 fanout648 (.A(net649),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net652),
    .X(net649));
 sg13g2_buf_8 fanout650 (.A(net652),
    .X(net650));
 sg13g2_buf_8 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(net658),
    .X(net652));
 sg13g2_buf_8 fanout653 (.A(net657),
    .X(net653));
 sg13g2_buf_8 fanout654 (.A(net657),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_8 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_8 fanout658 (.A(net701),
    .X(net658));
 sg13g2_buf_8 fanout659 (.A(net661),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_8 fanout661 (.A(net664),
    .X(net661));
 sg13g2_buf_8 fanout662 (.A(net664),
    .X(net662));
 sg13g2_buf_8 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_8 fanout664 (.A(net667),
    .X(net664));
 sg13g2_buf_8 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_8 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_8 fanout667 (.A(net701),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(net671),
    .X(net668));
 sg13g2_buf_8 fanout669 (.A(net671),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_8 fanout671 (.A(net675),
    .X(net671));
 sg13g2_buf_8 fanout672 (.A(net675),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(net675),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_8 fanout675 (.A(net701),
    .X(net675));
 sg13g2_buf_8 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_8 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_8 fanout678 (.A(net690),
    .X(net678));
 sg13g2_buf_8 fanout679 (.A(net682),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net682),
    .X(net680));
 sg13g2_buf_8 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_8 fanout682 (.A(net690),
    .X(net682));
 sg13g2_buf_8 fanout683 (.A(net685),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(net690),
    .X(net685));
 sg13g2_buf_8 fanout686 (.A(net689),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_8 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_8 fanout690 (.A(net701),
    .X(net690));
 sg13g2_buf_8 fanout691 (.A(net700),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net700),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(net700),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(net697),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(net697),
    .X(net695));
 sg13g2_buf_8 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_8 fanout697 (.A(net700),
    .X(net697));
 sg13g2_buf_8 fanout698 (.A(net700),
    .X(net698));
 sg13g2_buf_8 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_8 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_8 fanout701 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.rstn ),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(_0954_),
    .X(net702));
 sg13g2_buf_8 fanout703 (.A(_0449_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_0449_),
    .X(net704));
 sg13g2_buf_8 fanout705 (.A(_2002_),
    .X(net705));
 sg13g2_buf_8 fanout706 (.A(_1986_),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(_1965_),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(_1963_),
    .X(net708));
 sg13g2_buf_8 fanout709 (.A(_1963_),
    .X(net709));
 sg13g2_buf_8 fanout710 (.A(net712),
    .X(net710));
 sg13g2_buf_1 fanout711 (.A(net713),
    .X(net711));
 sg13g2_buf_8 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_8 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(_1929_),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(_1916_),
    .X(net715));
 sg13g2_buf_1 fanout716 (.A(_1916_),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(_1900_),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(_1897_),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(_1896_),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(_1895_),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(_1894_),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(net724),
    .X(net722));
 sg13g2_buf_8 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(net733),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(net733),
    .X(net726));
 sg13g2_buf_8 fanout727 (.A(net733),
    .X(net727));
 sg13g2_buf_8 fanout728 (.A(net732),
    .X(net728));
 sg13g2_buf_8 fanout729 (.A(net732),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_8 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_8 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_8 fanout733 (.A(net734),
    .X(net733));
 sg13g2_buf_8 fanout734 (.A(net1036),
    .X(net734));
 sg13g2_buf_8 fanout735 (.A(net737),
    .X(net735));
 sg13g2_buf_8 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_8 fanout737 (.A(\u_usb_cdc.clk_gate_q ),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_8 fanout739 (.A(net744),
    .X(net739));
 sg13g2_buf_8 fanout740 (.A(net742),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_8 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_8 fanout743 (.A(net744),
    .X(net743));
 sg13g2_buf_8 fanout744 (.A(net1049),
    .X(net744));
 sg13g2_buf_8 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_8 fanout746 (.A(net976),
    .X(net746));
 sg13g2_buf_8 fanout747 (.A(net944),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net944),
    .X(net748));
 sg13g2_buf_8 fanout749 (.A(net1068),
    .X(net749));
 sg13g2_buf_8 fanout750 (.A(net1044),
    .X(net750));
 sg13g2_buf_8 fanout751 (.A(net942),
    .X(net751));
 sg13g2_buf_8 fanout752 (.A(net991),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net1014),
    .X(net753));
 sg13g2_buf_8 fanout754 (.A(net996),
    .X(net754));
 sg13g2_buf_8 fanout755 (.A(net1016),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(net1062),
    .X(net756));
 sg13g2_buf_8 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_8 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_8 fanout759 (.A(\u_usb_cdc.sie_out_data[1] ),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_8 fanout761 (.A(net399),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(net763),
    .X(net762));
 sg13g2_buf_8 fanout763 (.A(net1023),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_8 fanout765 (.A(net1052),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(net986),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(\u_usb_cdc.endp[0] ),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net1056),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(net772),
    .X(net770));
 sg13g2_buf_1 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(net1031),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(net775),
    .X(net773));
 sg13g2_buf_1 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_8 fanout775 (.A(net1030),
    .X(net775));
 sg13g2_buf_8 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_8 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(net1061),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net782),
    .X(net780));
 sg13g2_buf_1 fanout781 (.A(net782),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(net1060),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(net1043),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_8 fanout787 (.A(net1063),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net1048),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net790),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net796),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(net796),
    .X(net794));
 sg13g2_buf_1 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(net1026),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net804),
    .X(net797));
 sg13g2_buf_8 fanout798 (.A(net804),
    .X(net798));
 sg13g2_buf_8 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_8 fanout800 (.A(net804),
    .X(net800));
 sg13g2_buf_8 fanout801 (.A(net802),
    .X(net801));
 sg13g2_buf_8 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[0] ),
    .X(net804));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805));
 sg13g2_buf_8 fanout806 (.A(net1064),
    .X(net806));
 sg13g2_buf_8 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_8 fanout808 (.A(net1024),
    .X(net808));
 sg13g2_buf_8 fanout809 (.A(net810),
    .X(net809));
 sg13g2_buf_8 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_8 fanout811 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[1] ),
    .X(net811));
 sg13g2_buf_8 fanout812 (.A(net814),
    .X(net812));
 sg13g2_buf_1 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_8 fanout814 (.A(net819),
    .X(net814));
 sg13g2_buf_8 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_8 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_8 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_8 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_8 fanout819 (.A(net1054),
    .X(net819));
 sg13g2_buf_8 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_8 fanout821 (.A(net1057),
    .X(net821));
 sg13g2_buf_8 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_8 fanout823 (.A(net1059),
    .X(net823));
 sg13g2_buf_8 fanout824 (.A(net826),
    .X(net824));
 sg13g2_buf_1 fanout825 (.A(net826),
    .X(net825));
 sg13g2_buf_8 fanout826 (.A(net1065),
    .X(net826));
 sg13g2_buf_8 fanout827 (.A(net1053),
    .X(net827));
 sg13g2_buf_8 fanout828 (.A(net1067),
    .X(net828));
 sg13g2_buf_8 fanout829 (.A(net561),
    .X(net829));
 sg13g2_buf_8 fanout830 (.A(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .X(net830));
 sg13g2_buf_8 fanout831 (.A(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .X(net831));
 sg13g2_buf_8 fanout832 (.A(net981),
    .X(net832));
 sg13g2_buf_8 fanout833 (.A(net847),
    .X(net833));
 sg13g2_buf_8 fanout834 (.A(net835),
    .X(net834));
 sg13g2_buf_8 fanout835 (.A(net1045),
    .X(net835));
 sg13g2_buf_8 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_8 fanout837 (.A(\u_usb_cdc.u_sie.phy_state_q[6] ),
    .X(net837));
 sg13g2_buf_8 fanout838 (.A(net939),
    .X(net838));
 sg13g2_buf_8 fanout839 (.A(\u_usb_cdc.u_sie.phy_state_q[1] ),
    .X(net839));
 sg13g2_buf_1 fanout840 (.A(net1050),
    .X(net840));
 sg13g2_buf_8 fanout841 (.A(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .X(net841));
 sg13g2_buf_8 fanout842 (.A(net1029),
    .X(net842));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(usb_dn_rx_i),
    .X(net12));
 sg13g2_buf_1 input13 (.A(usb_dp_rx_i),
    .X(net13));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[2]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[3]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[4]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[5]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[6]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_oe[7]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[0]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[1]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[2]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[3]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[4]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[5]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uio_out[6]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[0]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[1]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[2]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[3]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[4]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[5]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[6]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(uo_out[7]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(usb_dn_en_o));
 sg13g2_buf_1 output38 (.A(net38),
    .X(usb_dn_tx_o));
 sg13g2_buf_1 output39 (.A(net39),
    .X(usb_dp_en_o));
 sg13g2_buf_1 output40 (.A(net40),
    .X(usb_dp_tx_o));
 sg13g2_tielo heichips25_usb_cdc_41 (.L_LO(net41));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload0 (.A(clknet_leaf_55_clk));
 sg13g2_inv_4 clkload1 (.A(clknet_leaf_48_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_leaf_35_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_29_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_usb_cdc.u_sie.u_phy_rx.dn_q[2] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_usb_cdc.u_sie.u_phy_rx.dp_q[2] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_usb_cdc.rstn_sq[1] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_usb_cdc.u_sie.u_phy_rx.dn_q[1] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_usb_cdc.u_sie.u_phy_rx.dp_q[1] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_usb_cdc.clk_cnt_q[0] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[0] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0046_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_usb_cdc.clk_cnt_q[1] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[2] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0401_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[6] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0173_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[45] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0128_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[27] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[55] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0138_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[20] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0103_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[3] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold22 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[44] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0211_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[26] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[23] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0106_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[12] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0095_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[46] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0129_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[41] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0124_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[9] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0092_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[35] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[40] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0207_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[47] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0130_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[2] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[40] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0123_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_usb_cdc.u_sie.in_zlp_q[1] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0436_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[54] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0137_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[17] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0100_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[15] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0098_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[21] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0104_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[8] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0091_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[1] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[37] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0204_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[68] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0235_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[11] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0178_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[8] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0175_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[53] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0136_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[45] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0212_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[42] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0125_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[47] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0214_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[49] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0132_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold74 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[70] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0237_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[64] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0231_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[66] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0233_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[10] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0177_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[50] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0133_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[52] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0135_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[62] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0229_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[44] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0127_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold90 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[42] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0209_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[69] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0236_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0052_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[11] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0094_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[38] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0205_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold99 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[39] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0206_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold101 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[71] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0238_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold103 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[65] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0232_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold105 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[22] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0105_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold107 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[43] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0126_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[14] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0097_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[12] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0179_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[48] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0131_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold115 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[4] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0171_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[51] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0134_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[63] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[16] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0099_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[59] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_usb_cdc.u_sie.in_zlp_q[0] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0437_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[61] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0228_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_usb_cdc.u_sie.out_toggle_q[0] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0989_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0067_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[6] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0387_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[34] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold133 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[58] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold134 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[28] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0195_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[18] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0101_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold138 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[14] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0181_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold140 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[30] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0197_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold142 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[19] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0102_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_usb_cdc.u_sie.phy_state_q[5] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0024_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[33] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[17] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0398_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold149 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[10] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0093_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold151 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[67] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0234_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[43] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0210_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[46] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0213_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[57] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold158 (.A(\u_usb_cdc.u_sie.addr_q[3] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[31] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[2] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0383_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[29] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0196_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold164 (.A(\u_usb_cdc.u_ctrl_endp.req_q[10] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0000_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0050_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0025_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0058_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[2] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0423_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold171 (.A(\u_usb_cdc.u_sie.addr_q[2] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_usb_cdc.u_sie.addr_q[5] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0311_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[9] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0176_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_usb_cdc.u_sie.addr_q[0] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold177 (.A(_1030_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0072_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[15] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0182_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[56] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0223_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[13] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0180_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[24] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0191_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[7] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold188 (.A(\u_usb_cdc.u_sie.in_byte_q[2] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0321_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold190 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[5] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0172_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_usb_cdc.dp_pu_o ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold193 (.A(_1804_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0420_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_usb_cdc.u_sie.addr_q[4] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0310_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[25] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold198 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[36] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0203_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold200 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[32] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0199_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold202 (.A(\u_usb_cdc.u_sie.u_phy_rx.se0_q ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0432_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold204 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[41] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0208_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold206 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[60] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0227_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_usb_cdc.u_sie.addr_q[6] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0312_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_usb_cdc.u_sie.addr_q[1] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[13] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0096_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[0] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0167_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold215 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[4] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0032_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold217 (.A(\u_usb_cdc.u_sie.phy_state_q[10] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0584_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0596_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0063_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold221 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_err_q ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0974_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[3] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0424_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold225 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[22] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0189_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold227 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[0] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0268_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold229 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[3] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold230 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[55] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0222_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[5] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0426_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold234 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[50] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0217_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold236 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[4] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0385_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold238 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[2] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0165_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold240 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[1] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[21] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0188_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold243 (.A(\u_usb_cdc.u_sie.crc16_q[4] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0335_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold245 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[5] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0386_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold247 (.A(\u_usb_cdc.u_sie.in_byte_q[0] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0319_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_usb_cdc.u_sie.out_eop_q ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold250 (.A(_1717_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0371_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold252 (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[1] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold253 (.A(_1792_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0400_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold255 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[14] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0395_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold257 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[20] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0187_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold259 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[0] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0163_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold261 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[10] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0391_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold263 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[15] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold264 (.A(\u_usb_cdc.u_sie.crc16_q[5] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0336_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0054_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0073_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_usb_cdc.u_sie.in_toggle_q[0] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0069_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0059_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0430_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold272 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[23] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0190_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold274 (.A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[1] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0434_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold276 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[0] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold277 (.A(\u_usb_cdc.u_sie.in_byte_q[1] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0320_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold279 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[18] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0185_),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold281 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[52] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0219_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold283 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[51] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0218_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold285 (.A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[0] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0433_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold287 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[54] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0221_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold289 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0382_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold291 (.A(\u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q[2] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0435_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold293 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[3] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0166_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[63] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0146_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold297 (.A(\u_usb_cdc.u_sie.in_byte_q[3] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0322_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold299 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[2] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold300 (.A(\u_usb_cdc.u_sie.u_phy_rx.state_q[1] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0950_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0033_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold303 (.A(\u_usb_cdc.u_ctrl_endp.dev_state_q[1] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold304 (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[1] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold305 (.A(_1461_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0314_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold307 (.A(\u_usb_cdc.u_sie.crc16_q[6] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0337_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0051_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0456_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0064_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold312 (.A(\u_usb_cdc.u_sie.in_toggle_q[2] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1025_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0071_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold315 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold316 (.A(_1796_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0403_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0056_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0419_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold320 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[48] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0215_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold322 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[6] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0281_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold324 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[13] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0394_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0057_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0428_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold328 (.A(net19),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0360_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold330 (.A(\u_usb_cdc.u_sie.crc16_q[3] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0334_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold332 (.A(net16),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0357_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold334 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[39] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0122_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold336 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[0] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0083_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold338 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[6] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0089_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0053_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0037_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold342 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[4] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0279_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold344 (.A(\u_usb_cdc.u_sie.u_phy_rx.dn_q[0] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold345 (.A(_1802_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0410_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold347 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[16] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0183_),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold349 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[1] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold351 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[9] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0390_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold353 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[56] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0139_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold355 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[4] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0087_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold357 (.A(\u_usb_cdc.sie_out_data[0] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold358 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[6] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold359 (.A(_1862_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold360 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[8] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0389_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold362 (.A(net29),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold363 (.A(_1276_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0243_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold365 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[3] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0086_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold367 (.A(\u_usb_cdc.u_sie.crc16_q[0] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold368 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[29] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0112_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold370 (.A(net14),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold371 (.A(\u_usb_cdc.u_sie.phy_state_q[2] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0021_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0055_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold374 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[49] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0216_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold376 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[24] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0107_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold378 (.A(net15),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0356_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold380 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[11] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold381 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[1] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold382 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0085_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold384 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[26] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0109_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold386 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[5] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold387 (.A(_1725_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold388 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[65] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0148_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold390 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[69] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0152_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold392 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[57] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0140_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold394 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[32] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0115_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold396 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[7] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0090_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold398 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[19] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0186_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold400 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[1] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0084_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold402 (.A(\u_usb_cdc.u_sie.crc16_q[10] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0523_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold404 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[34] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0117_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold406 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[68] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0151_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold408 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[64] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0147_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold410 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[27] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0110_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold412 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[35] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0118_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold414 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[30] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0113_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold416 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[5] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0280_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold418 (.A(\u_usb_cdc.u_sie.delay_cnt_q[2] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0318_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold420 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[62] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0145_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold422 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[66] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0149_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold424 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[4] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold425 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[36] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0119_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold427 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[70] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0153_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold429 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[33] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0116_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold431 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[31] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0114_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold433 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[38] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0121_),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold435 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[67] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0150_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold437 (.A(\u_usb_cdc.u_ctrl_endp.in_endp_q ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0267_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold439 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[28] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0111_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold441 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[61] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0144_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold443 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[2] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold444 (.A(_1722_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold445 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[60] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0143_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold447 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[25] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0108_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold449 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[71] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0154_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold451 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[59] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0142_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold453 (.A(net31),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0245_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold455 (.A(\u_usb_cdc.u_sie.u_phy_rx.state_q[2] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0951_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold457 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[53] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold458 (.A(_1217_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0220_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold460 (.A(\u_usb_cdc.u_sie.crc16_q[2] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold461 (.A(net20),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0361_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold463 (.A(net17),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0358_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold465 (.A(\u_usb_cdc.u_sie.delay_cnt_q[1] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold466 (.A(_1470_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0317_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold468 (.A(\u_usb_cdc.u_ctrl_endp.addr_dd[3] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold469 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[58] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0141_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold471 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[37] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0120_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold473 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[3] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold474 (.A(_1735_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0380_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold476 (.A(\u_usb_cdc.u_ctrl_endp.endp_q[0] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold477 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_eop_q ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0975_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold479 (.A(\u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q[1] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0047_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold481 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[2] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0290_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold483 (.A(\u_usb_cdc.u_sie.phy_state_q[3] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0022_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold485 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[4] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold486 (.A(_1724_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold487 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_valid_q ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0045_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold489 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[1] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold490 (.A(_1721_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold491 (.A(\u_usb_cdc.out_valid_o [0]),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0042_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0049_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0642_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0062_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold496 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[4] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0292_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold498 (.A(\u_usb_cdc.u_sie.crc16_q[9] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0501_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold500 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0074_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold502 (.A(net33),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0247_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold504 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_fifo_q[17] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0184_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold506 (.A(\u_usb_cdc.u_sie.crc16_q[12] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0518_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold508 (.A(\u_usb_cdc.u_ctrl_endp.state_q[1] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0011_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold510 (.A(\u_usb_cdc.u_ctrl_endp.req_q[11] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0001_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold512 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_fifo_q[5] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0088_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold514 (.A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[1] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold515 (.A(_0955_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0036_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold517 (.A(net32),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0246_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold519 (.A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[3] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0958_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold521 (.A(\u_usb_cdc.u_sie.crc16_q[13] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold522 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold523 (.A(_1892_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold524 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[16] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold525 (.A(net21),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0362_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold527 (.A(\u_usb_cdc.u_ctrl_endp.req_q[8] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0009_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold529 (.A(\u_usb_cdc.u_sie.phy_state_q[8] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0027_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold531 (.A(\u_usb_cdc.u_sie.out_toggle_q[1] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold532 (.A(_1002_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0068_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold534 (.A(\u_usb_cdc.u_sie.u_phy_rx.dp_q[0] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold535 (.A(_0409_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold536 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[5] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0293_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold538 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[1] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold539 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[2] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold540 (.A(net18),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold541 (.A(_0359_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0048_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0061_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold544 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[6] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold545 (.A(_1726_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold546 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[0] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold547 (.A(\u_usb_cdc.addr[5] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold548 (.A(\u_usb_cdc.u_ctrl_endp.state_q[5] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0015_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold550 (.A(\u_usb_cdc.u_ctrl_endp.req_q[1] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0002_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold552 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[1] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold553 (.A(\u_usb_cdc.u_ctrl_endp.state_q[3] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0013_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold555 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[7] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold556 (.A(net36),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold557 (.A(_0250_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold558 (.A(net35),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0249_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold560 (.A(\u_usb_cdc.bus_reset ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0402_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold562 (.A(\u_usb_cdc.addr[1] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold563 (.A(\u_usb_cdc.u_sie.crc16_q[8] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold564 (.A(\u_usb_cdc.u_sie.crc16_q[7] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0330_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold566 (.A(\u_usb_cdc.u_ctrl_endp.class_q ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold567 (.A(_0286_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold568 (.A(\u_usb_cdc.addr[6] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[12] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold570 (.A(\u_usb_cdc.u_ctrl_endp.state_q[7] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0017_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold572 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[6] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0294_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold574 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[1] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0029_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold576 (.A(net30),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0244_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold578 (.A(\u_usb_cdc.addr[4] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold579 (.A(net34),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0248_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold581 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[3] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold582 (.A(_1723_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold583 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[3] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold584 (.A(_0157_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold585 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_qq[0] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold586 (.A(\u_usb_cdc.u_sie.pid_q[0] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold587 (.A(\u_usb_cdc.addr[3] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold588 (.A(\u_usb_cdc.u_ctrl_endp.req_q[6] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0007_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold590 (.A(\u_usb_cdc.u_sie.u_phy_rx.shift_register_q[7] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold591 (.A(_1727_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold592 (.A(\u_usb_cdc.u_ctrl_endp.rec_q[1] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold593 (.A(net26),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0363_),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold595 (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[1] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0408_),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold597 (.A(\u_usb_cdc.u_sie.crc16_q[15] ),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold598 (.A(\u_usb_cdc.u_ctrl_endp.max_length_q[3] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold599 (.A(_0291_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold600 (.A(\u_usb_cdc.u_sie.crc16_q[1] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold601 (.A(\u_usb_cdc.u_sie.data_q[7] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold602 (.A(\u_usb_cdc.u_ctrl_endp.rec_q[0] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold603 (.A(\u_usb_cdc.u_ctrl_endp.req_q[7] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0008_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold605 (.A(\u_usb_cdc.u_sie.in_toggle_q[1] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold606 (.A(_1021_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold607 (.A(_0070_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold608 (.A(\u_usb_cdc.addr[2] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold609 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_q[1] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold610 (.A(_0164_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold611 (.A(\u_usb_cdc.u_sie.rx_data[4] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0416_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold613 (.A(\u_usb_cdc.u_sie.u_phy_tx.tx_state_q[2] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold614 (.A(_0066_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold615 (.A(net28),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0365_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold617 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_en_q ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold618 (.A(_0405_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold619 (.A(\u_usb_cdc.u_ctrl_endp.dev_state_qq[0] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold620 (.A(_0313_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold621 (.A(\u_usb_cdc.u_sie.phy_state_q[4] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold622 (.A(\u_usb_cdc.u_sie.rx_data[1] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold623 (.A(\u_usb_cdc.in_ready_o [0]),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold624 (.A(\u_usb_cdc.sie_out_data[7] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold625 (.A(_0303_),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold626 (.A(\u_usb_cdc.u_sie.rx_err ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold627 (.A(\u_usb_cdc.u_sie.rx_data[2] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold628 (.A(\u_usb_cdc.ctrl_stall ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold629 (.A(_0859_),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0014_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold631 (.A(\u_usb_cdc.u_ctrl_endp.req_q[9] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold632 (.A(_0010_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold633 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[6] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold634 (.A(_0301_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold635 (.A(\u_usb_cdc.u_ctrl_endp.req_q[3] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold636 (.A(_0004_),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold637 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[0] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold638 (.A(_0251_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold639 (.A(\u_usb_cdc.u_sie.pid_q[1] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold640 (.A(\u_usb_cdc.endp[1] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0304_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold642 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[3] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold643 (.A(_0254_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold644 (.A(net27),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold645 (.A(_0364_),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold646 (.A(\u_usb_cdc.endp[3] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold647 (.A(_0306_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold648 (.A(\u_usb_cdc.u_sie.rx_data[3] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold649 (.A(\u_usb_cdc.u_sie.rx_data[0] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold650 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[1] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold651 (.A(_0252_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold652 (.A(\u_usb_cdc.u_ctrl_endp.req_q[2] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold653 (.A(\u_usb_cdc.u_ctrl_endp.req_q[4] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold654 (.A(_0005_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold655 (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[0] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold656 (.A(_0407_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold657 (.A(\u_usb_cdc.u_sie.phy_state_q[11] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold658 (.A(\u_usb_cdc.u_sie.rx_valid ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold659 (.A(_1800_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold660 (.A(_0406_),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold661 (.A(\u_usb_cdc.u_sie.u_phy_tx.data_q[0] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold662 (.A(\u_usb_cdc.u_sie.data_q[4] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold663 (.A(\u_usb_cdc.u_sie.phy_state_q[9] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold664 (.A(\u_usb_cdc.u_sie.rx_data[6] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold665 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_q[2] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold666 (.A(_0253_),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold667 (.A(\u_usb_cdc.u_sie.data_q[6] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold668 (.A(\u_usb_cdc.u_sie.data_q[0] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold669 (.A(\u_usb_cdc.u_sie.u_phy_rx.state_q[3] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold670 (.A(\u_usb_cdc.u_sie.u_phy_rx.nrzi_q[2] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold671 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[2] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold672 (.A(_0261_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold673 (.A(\u_usb_cdc.sie_out_data[6] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold674 (.A(\u_usb_cdc.u_sie.rx_data[5] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold675 (.A(\u_usb_cdc.u_ctrl_endp.in_dir_q ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold676 (.A(\u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q[0] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold677 (.A(\u_usb_cdc.u_sie.data_q[5] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold678 (.A(\u_usb_cdc.sie_out_data[4] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold679 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0159_),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold681 (.A(\u_usb_cdc.u_sie.rx_data[7] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold682 (.A(_0060_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold683 (.A(_1873_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold684 (.A(\u_usb_cdc.endp[2] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold685 (.A(\u_usb_cdc.u_ctrl_endp.state_q[6] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold686 (.A(_0016_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold687 (.A(\u_usb_cdc.u_sie.delay_cnt_q[0] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold688 (.A(_0316_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold689 (.A(\u_usb_cdc.u_sie.u_phy_rx.cnt_q[3] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold690 (.A(_0384_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold691 (.A(\u_usb_cdc.u_sie.pid_q[2] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold692 (.A(_0368_),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold693 (.A(\u_usb_cdc.u_sie.data_q[3] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold694 (.A(\u_usb_cdc.u_sie.u_phy_rx.rx_state_q[2] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold695 (.A(_0030_),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold696 (.A(\u_usb_cdc.sie_out_data[5] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold697 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[1] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold698 (.A(\u_usb_cdc.sie_out_data[3] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold699 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold700 (.A(\u_usb_cdc.u_sie.pid_q[3] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold701 (.A(_0369_),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold702 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[3] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold703 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[1] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold704 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[0] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold705 (.A(\u_usb_cdc.u_sie.data_q[2] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold706 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[2] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold707 (.A(_0257_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold708 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[1] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold709 (.A(_1367_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold710 (.A(_0260_),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold711 (.A(\u_usb_cdc.u_ctrl_endp.req_q[5] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold712 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[4] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold713 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[5] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold714 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[2] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold715 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[4] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold716 (.A(\u_usb_cdc.sie_in_data_ack ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold717 (.A(_0411_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold718 (.A(\u_usb_cdc.rstn ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold719 (.A(\u_usb_cdc.u_ctrl_endp.state_q[2] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold720 (.A(_0855_),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold721 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[7] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold722 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[3] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold723 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[5] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold724 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q[6] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold725 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[1] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold726 (.A(\u_usb_cdc.sie_out_err ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold727 (.A(\u_usb_cdc.u_sie.phy_state_q[7] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold728 (.A(\u_usb_cdc.sie_in_req ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold729 (.A(_0259_),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold730 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_first_qq[3] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold731 (.A(\u_usb_cdc.clk_gate_q ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold732 (.A(\u_usb_cdc.u_sie.phy_state_q[1] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold733 (.A(_0020_),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold734 (.A(\u_usb_cdc.u_sie.data_q[1] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold735 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold736 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[0] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold737 (.A(_0255_),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold738 (.A(\u_usb_cdc.bulk_out_nak [0]),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold739 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[2] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold740 (.A(_0241_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold741 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[0] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold742 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[2] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold743 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[3] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold744 (.A(\u_usb_cdc.sie_out_data[2] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold745 (.A(\u_usb_cdc.u_ctrl_endp.byte_cnt_q[0] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold746 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_first_q[3] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold747 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[2] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold748 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[1] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold749 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_in_fifo.in_last_q[0] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold750 (.A(\u_usb_cdc.sie_out_err ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold751 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold752 (.A(\u_usb_cdc.u_bulk_endps[0].u_bulk_endp.u_out_fifo.out_last_qq[3] ),
    .X(net1070));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_56 ();
 sg13g2_fill_1 FILLER_0_89 ();
 sg13g2_decap_4 FILLER_0_107 ();
 sg13g2_fill_1 FILLER_0_111 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_fill_2 FILLER_0_133 ();
 sg13g2_fill_2 FILLER_0_153 ();
 sg13g2_decap_4 FILLER_0_209 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_fill_2 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_fill_2 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_0_409 ();
 sg13g2_decap_8 FILLER_0_416 ();
 sg13g2_decap_8 FILLER_0_423 ();
 sg13g2_decap_8 FILLER_0_430 ();
 sg13g2_decap_8 FILLER_0_437 ();
 sg13g2_decap_8 FILLER_0_444 ();
 sg13g2_decap_8 FILLER_0_451 ();
 sg13g2_decap_8 FILLER_0_458 ();
 sg13g2_decap_8 FILLER_0_465 ();
 sg13g2_decap_8 FILLER_0_472 ();
 sg13g2_decap_8 FILLER_0_479 ();
 sg13g2_decap_8 FILLER_0_486 ();
 sg13g2_decap_8 FILLER_0_493 ();
 sg13g2_decap_8 FILLER_0_500 ();
 sg13g2_decap_8 FILLER_0_507 ();
 sg13g2_decap_8 FILLER_0_514 ();
 sg13g2_decap_8 FILLER_0_521 ();
 sg13g2_decap_8 FILLER_0_528 ();
 sg13g2_decap_8 FILLER_0_535 ();
 sg13g2_decap_8 FILLER_0_542 ();
 sg13g2_decap_8 FILLER_0_549 ();
 sg13g2_decap_8 FILLER_0_556 ();
 sg13g2_decap_8 FILLER_0_563 ();
 sg13g2_decap_8 FILLER_0_570 ();
 sg13g2_decap_8 FILLER_0_577 ();
 sg13g2_decap_8 FILLER_0_584 ();
 sg13g2_decap_8 FILLER_0_591 ();
 sg13g2_decap_8 FILLER_0_598 ();
 sg13g2_decap_8 FILLER_0_605 ();
 sg13g2_decap_8 FILLER_0_612 ();
 sg13g2_decap_8 FILLER_0_619 ();
 sg13g2_decap_8 FILLER_0_626 ();
 sg13g2_decap_8 FILLER_0_633 ();
 sg13g2_decap_8 FILLER_0_640 ();
 sg13g2_decap_8 FILLER_0_647 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_8 FILLER_0_661 ();
 sg13g2_decap_8 FILLER_0_668 ();
 sg13g2_decap_8 FILLER_0_675 ();
 sg13g2_decap_8 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_4 FILLER_0_1025 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_fill_2 FILLER_1_21 ();
 sg13g2_fill_2 FILLER_1_37 ();
 sg13g2_fill_1 FILLER_1_74 ();
 sg13g2_fill_1 FILLER_1_111 ();
 sg13g2_fill_1 FILLER_1_166 ();
 sg13g2_fill_2 FILLER_1_199 ();
 sg13g2_fill_1 FILLER_1_201 ();
 sg13g2_decap_4 FILLER_1_265 ();
 sg13g2_fill_1 FILLER_1_269 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_fill_2 FILLER_1_281 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_decap_8 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_1_435 ();
 sg13g2_decap_8 FILLER_1_442 ();
 sg13g2_decap_8 FILLER_1_449 ();
 sg13g2_decap_8 FILLER_1_456 ();
 sg13g2_decap_8 FILLER_1_463 ();
 sg13g2_decap_8 FILLER_1_470 ();
 sg13g2_decap_8 FILLER_1_477 ();
 sg13g2_decap_8 FILLER_1_484 ();
 sg13g2_decap_8 FILLER_1_491 ();
 sg13g2_decap_8 FILLER_1_498 ();
 sg13g2_decap_8 FILLER_1_505 ();
 sg13g2_decap_8 FILLER_1_512 ();
 sg13g2_decap_8 FILLER_1_519 ();
 sg13g2_decap_8 FILLER_1_526 ();
 sg13g2_decap_8 FILLER_1_533 ();
 sg13g2_decap_8 FILLER_1_540 ();
 sg13g2_decap_8 FILLER_1_547 ();
 sg13g2_decap_8 FILLER_1_554 ();
 sg13g2_decap_8 FILLER_1_561 ();
 sg13g2_decap_8 FILLER_1_568 ();
 sg13g2_decap_8 FILLER_1_575 ();
 sg13g2_decap_8 FILLER_1_582 ();
 sg13g2_decap_8 FILLER_1_589 ();
 sg13g2_decap_8 FILLER_1_596 ();
 sg13g2_decap_8 FILLER_1_603 ();
 sg13g2_decap_8 FILLER_1_610 ();
 sg13g2_decap_8 FILLER_1_617 ();
 sg13g2_decap_8 FILLER_1_624 ();
 sg13g2_decap_8 FILLER_1_631 ();
 sg13g2_decap_8 FILLER_1_638 ();
 sg13g2_decap_8 FILLER_1_645 ();
 sg13g2_decap_8 FILLER_1_652 ();
 sg13g2_decap_8 FILLER_1_659 ();
 sg13g2_decap_8 FILLER_1_666 ();
 sg13g2_decap_8 FILLER_1_673 ();
 sg13g2_decap_8 FILLER_1_680 ();
 sg13g2_decap_8 FILLER_1_687 ();
 sg13g2_decap_8 FILLER_1_694 ();
 sg13g2_decap_8 FILLER_1_701 ();
 sg13g2_decap_8 FILLER_1_708 ();
 sg13g2_decap_8 FILLER_1_715 ();
 sg13g2_decap_8 FILLER_1_722 ();
 sg13g2_decap_8 FILLER_1_729 ();
 sg13g2_decap_8 FILLER_1_736 ();
 sg13g2_decap_8 FILLER_1_743 ();
 sg13g2_decap_8 FILLER_1_750 ();
 sg13g2_decap_8 FILLER_1_757 ();
 sg13g2_decap_8 FILLER_1_764 ();
 sg13g2_decap_8 FILLER_1_771 ();
 sg13g2_decap_8 FILLER_1_778 ();
 sg13g2_decap_8 FILLER_1_785 ();
 sg13g2_decap_8 FILLER_1_792 ();
 sg13g2_decap_8 FILLER_1_799 ();
 sg13g2_decap_8 FILLER_1_806 ();
 sg13g2_decap_8 FILLER_1_813 ();
 sg13g2_decap_8 FILLER_1_820 ();
 sg13g2_decap_8 FILLER_1_827 ();
 sg13g2_decap_8 FILLER_1_834 ();
 sg13g2_decap_8 FILLER_1_841 ();
 sg13g2_decap_8 FILLER_1_848 ();
 sg13g2_decap_8 FILLER_1_855 ();
 sg13g2_decap_8 FILLER_1_862 ();
 sg13g2_decap_8 FILLER_1_869 ();
 sg13g2_decap_8 FILLER_1_876 ();
 sg13g2_decap_8 FILLER_1_883 ();
 sg13g2_decap_8 FILLER_1_890 ();
 sg13g2_decap_8 FILLER_1_897 ();
 sg13g2_decap_8 FILLER_1_904 ();
 sg13g2_decap_8 FILLER_1_911 ();
 sg13g2_decap_8 FILLER_1_918 ();
 sg13g2_decap_8 FILLER_1_925 ();
 sg13g2_decap_8 FILLER_1_932 ();
 sg13g2_decap_8 FILLER_1_939 ();
 sg13g2_decap_8 FILLER_1_946 ();
 sg13g2_decap_8 FILLER_1_953 ();
 sg13g2_decap_8 FILLER_1_960 ();
 sg13g2_decap_8 FILLER_1_967 ();
 sg13g2_decap_8 FILLER_1_974 ();
 sg13g2_decap_8 FILLER_1_981 ();
 sg13g2_decap_8 FILLER_1_988 ();
 sg13g2_decap_8 FILLER_1_995 ();
 sg13g2_decap_8 FILLER_1_1002 ();
 sg13g2_decap_8 FILLER_1_1009 ();
 sg13g2_decap_8 FILLER_1_1016 ();
 sg13g2_decap_4 FILLER_1_1023 ();
 sg13g2_fill_2 FILLER_1_1027 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_fill_1 FILLER_2_11 ();
 sg13g2_fill_1 FILLER_2_48 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_4 FILLER_2_105 ();
 sg13g2_fill_1 FILLER_2_109 ();
 sg13g2_fill_1 FILLER_2_155 ();
 sg13g2_decap_4 FILLER_2_205 ();
 sg13g2_fill_1 FILLER_2_209 ();
 sg13g2_decap_4 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_222 ();
 sg13g2_fill_2 FILLER_2_246 ();
 sg13g2_fill_1 FILLER_2_261 ();
 sg13g2_fill_2 FILLER_2_287 ();
 sg13g2_fill_2 FILLER_2_302 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_fill_2 FILLER_2_490 ();
 sg13g2_fill_1 FILLER_2_492 ();
 sg13g2_decap_4 FILLER_2_498 ();
 sg13g2_fill_2 FILLER_2_502 ();
 sg13g2_fill_2 FILLER_2_509 ();
 sg13g2_fill_1 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_516 ();
 sg13g2_fill_2 FILLER_2_523 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_8 ();
 sg13g2_decap_4 FILLER_3_15 ();
 sg13g2_decap_4 FILLER_3_47 ();
 sg13g2_fill_1 FILLER_3_51 ();
 sg13g2_fill_2 FILLER_3_66 ();
 sg13g2_fill_1 FILLER_3_68 ();
 sg13g2_fill_1 FILLER_3_92 ();
 sg13g2_fill_2 FILLER_3_103 ();
 sg13g2_decap_4 FILLER_3_132 ();
 sg13g2_fill_1 FILLER_3_163 ();
 sg13g2_decap_4 FILLER_3_195 ();
 sg13g2_fill_2 FILLER_3_203 ();
 sg13g2_fill_1 FILLER_3_205 ();
 sg13g2_decap_4 FILLER_3_220 ();
 sg13g2_fill_2 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_253 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_fill_2 FILLER_3_278 ();
 sg13g2_fill_1 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_286 ();
 sg13g2_decap_8 FILLER_3_293 ();
 sg13g2_fill_2 FILLER_3_313 ();
 sg13g2_fill_1 FILLER_3_315 ();
 sg13g2_fill_2 FILLER_3_321 ();
 sg13g2_decap_4 FILLER_3_337 ();
 sg13g2_fill_1 FILLER_3_341 ();
 sg13g2_fill_1 FILLER_3_351 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_fill_1 FILLER_3_391 ();
 sg13g2_fill_1 FILLER_3_397 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_4 FILLER_3_423 ();
 sg13g2_fill_1 FILLER_3_427 ();
 sg13g2_decap_4 FILLER_3_437 ();
 sg13g2_fill_2 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_452 ();
 sg13g2_decap_8 FILLER_3_459 ();
 sg13g2_decap_4 FILLER_3_466 ();
 sg13g2_fill_1 FILLER_3_470 ();
 sg13g2_fill_2 FILLER_3_534 ();
 sg13g2_decap_8 FILLER_3_545 ();
 sg13g2_fill_1 FILLER_3_552 ();
 sg13g2_decap_4 FILLER_3_562 ();
 sg13g2_fill_1 FILLER_3_566 ();
 sg13g2_decap_8 FILLER_3_572 ();
 sg13g2_decap_8 FILLER_3_579 ();
 sg13g2_decap_8 FILLER_3_586 ();
 sg13g2_decap_4 FILLER_3_593 ();
 sg13g2_fill_2 FILLER_3_597 ();
 sg13g2_decap_8 FILLER_3_626 ();
 sg13g2_decap_8 FILLER_3_633 ();
 sg13g2_decap_8 FILLER_3_640 ();
 sg13g2_decap_8 FILLER_3_647 ();
 sg13g2_decap_8 FILLER_3_654 ();
 sg13g2_decap_8 FILLER_3_661 ();
 sg13g2_decap_8 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_decap_8 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_689 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_decap_8 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_717 ();
 sg13g2_decap_8 FILLER_3_724 ();
 sg13g2_decap_8 FILLER_3_731 ();
 sg13g2_decap_8 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_745 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_3_878 ();
 sg13g2_decap_8 FILLER_3_885 ();
 sg13g2_decap_8 FILLER_3_892 ();
 sg13g2_decap_8 FILLER_3_899 ();
 sg13g2_decap_8 FILLER_3_906 ();
 sg13g2_decap_8 FILLER_3_913 ();
 sg13g2_decap_8 FILLER_3_920 ();
 sg13g2_decap_8 FILLER_3_927 ();
 sg13g2_decap_8 FILLER_3_934 ();
 sg13g2_decap_8 FILLER_3_941 ();
 sg13g2_decap_8 FILLER_3_948 ();
 sg13g2_decap_8 FILLER_3_955 ();
 sg13g2_decap_8 FILLER_3_962 ();
 sg13g2_decap_8 FILLER_3_969 ();
 sg13g2_decap_8 FILLER_3_976 ();
 sg13g2_decap_8 FILLER_3_983 ();
 sg13g2_decap_8 FILLER_3_990 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_4 FILLER_3_1025 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_2 FILLER_4_106 ();
 sg13g2_fill_1 FILLER_4_108 ();
 sg13g2_fill_1 FILLER_4_122 ();
 sg13g2_decap_8 FILLER_4_136 ();
 sg13g2_fill_2 FILLER_4_143 ();
 sg13g2_fill_1 FILLER_4_145 ();
 sg13g2_fill_1 FILLER_4_150 ();
 sg13g2_fill_2 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_273 ();
 sg13g2_fill_1 FILLER_4_296 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_4 FILLER_4_340 ();
 sg13g2_fill_2 FILLER_4_421 ();
 sg13g2_decap_8 FILLER_4_451 ();
 sg13g2_decap_8 FILLER_4_458 ();
 sg13g2_fill_1 FILLER_4_465 ();
 sg13g2_fill_2 FILLER_4_492 ();
 sg13g2_decap_8 FILLER_4_507 ();
 sg13g2_decap_8 FILLER_4_604 ();
 sg13g2_decap_8 FILLER_4_611 ();
 sg13g2_fill_1 FILLER_4_618 ();
 sg13g2_fill_1 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_641 ();
 sg13g2_decap_8 FILLER_4_648 ();
 sg13g2_decap_8 FILLER_4_655 ();
 sg13g2_decap_8 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_669 ();
 sg13g2_decap_8 FILLER_4_676 ();
 sg13g2_decap_8 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_decap_8 FILLER_4_704 ();
 sg13g2_decap_8 FILLER_4_711 ();
 sg13g2_decap_8 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_725 ();
 sg13g2_decap_8 FILLER_4_732 ();
 sg13g2_decap_8 FILLER_4_739 ();
 sg13g2_decap_8 FILLER_4_746 ();
 sg13g2_decap_8 FILLER_4_753 ();
 sg13g2_decap_8 FILLER_4_760 ();
 sg13g2_decap_8 FILLER_4_767 ();
 sg13g2_decap_8 FILLER_4_774 ();
 sg13g2_decap_8 FILLER_4_781 ();
 sg13g2_decap_8 FILLER_4_788 ();
 sg13g2_decap_8 FILLER_4_795 ();
 sg13g2_decap_8 FILLER_4_802 ();
 sg13g2_decap_8 FILLER_4_809 ();
 sg13g2_decap_8 FILLER_4_816 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_8 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_837 ();
 sg13g2_decap_8 FILLER_4_844 ();
 sg13g2_decap_8 FILLER_4_851 ();
 sg13g2_decap_8 FILLER_4_858 ();
 sg13g2_decap_8 FILLER_4_865 ();
 sg13g2_decap_8 FILLER_4_872 ();
 sg13g2_decap_8 FILLER_4_879 ();
 sg13g2_decap_8 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_893 ();
 sg13g2_decap_8 FILLER_4_900 ();
 sg13g2_decap_8 FILLER_4_907 ();
 sg13g2_decap_8 FILLER_4_914 ();
 sg13g2_decap_8 FILLER_4_921 ();
 sg13g2_decap_8 FILLER_4_928 ();
 sg13g2_decap_8 FILLER_4_935 ();
 sg13g2_decap_8 FILLER_4_942 ();
 sg13g2_decap_8 FILLER_4_949 ();
 sg13g2_decap_8 FILLER_4_956 ();
 sg13g2_decap_8 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_4 FILLER_4_1019 ();
 sg13g2_fill_2 FILLER_4_1023 ();
 sg13g2_fill_2 FILLER_5_4 ();
 sg13g2_fill_2 FILLER_5_52 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_decap_8 FILLER_5_72 ();
 sg13g2_decap_8 FILLER_5_79 ();
 sg13g2_fill_2 FILLER_5_86 ();
 sg13g2_fill_2 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_131 ();
 sg13g2_decap_8 FILLER_5_138 ();
 sg13g2_decap_4 FILLER_5_145 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_decap_4 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_222 ();
 sg13g2_fill_1 FILLER_5_224 ();
 sg13g2_decap_4 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_290 ();
 sg13g2_fill_2 FILLER_5_297 ();
 sg13g2_fill_2 FILLER_5_303 ();
 sg13g2_fill_2 FILLER_5_309 ();
 sg13g2_fill_1 FILLER_5_311 ();
 sg13g2_fill_1 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_4 FILLER_5_402 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_decap_4 FILLER_5_435 ();
 sg13g2_decap_8 FILLER_5_472 ();
 sg13g2_decap_8 FILLER_5_479 ();
 sg13g2_fill_1 FILLER_5_486 ();
 sg13g2_fill_2 FILLER_5_514 ();
 sg13g2_decap_8 FILLER_5_530 ();
 sg13g2_decap_4 FILLER_5_537 ();
 sg13g2_fill_2 FILLER_5_541 ();
 sg13g2_decap_8 FILLER_5_638 ();
 sg13g2_fill_2 FILLER_5_645 ();
 sg13g2_fill_1 FILLER_5_647 ();
 sg13g2_decap_8 FILLER_5_694 ();
 sg13g2_decap_8 FILLER_5_701 ();
 sg13g2_decap_8 FILLER_5_708 ();
 sg13g2_decap_8 FILLER_5_715 ();
 sg13g2_decap_8 FILLER_5_722 ();
 sg13g2_decap_8 FILLER_5_729 ();
 sg13g2_decap_8 FILLER_5_736 ();
 sg13g2_decap_8 FILLER_5_743 ();
 sg13g2_decap_8 FILLER_5_750 ();
 sg13g2_decap_8 FILLER_5_757 ();
 sg13g2_decap_8 FILLER_5_764 ();
 sg13g2_decap_8 FILLER_5_771 ();
 sg13g2_decap_8 FILLER_5_778 ();
 sg13g2_decap_8 FILLER_5_785 ();
 sg13g2_decap_8 FILLER_5_792 ();
 sg13g2_decap_8 FILLER_5_799 ();
 sg13g2_decap_8 FILLER_5_806 ();
 sg13g2_decap_8 FILLER_5_813 ();
 sg13g2_decap_8 FILLER_5_820 ();
 sg13g2_decap_8 FILLER_5_827 ();
 sg13g2_decap_8 FILLER_5_834 ();
 sg13g2_decap_8 FILLER_5_841 ();
 sg13g2_decap_8 FILLER_5_848 ();
 sg13g2_decap_8 FILLER_5_855 ();
 sg13g2_decap_8 FILLER_5_862 ();
 sg13g2_decap_8 FILLER_5_869 ();
 sg13g2_decap_8 FILLER_5_876 ();
 sg13g2_decap_8 FILLER_5_883 ();
 sg13g2_decap_8 FILLER_5_890 ();
 sg13g2_decap_8 FILLER_5_897 ();
 sg13g2_decap_8 FILLER_5_904 ();
 sg13g2_decap_8 FILLER_5_911 ();
 sg13g2_decap_8 FILLER_5_918 ();
 sg13g2_decap_8 FILLER_5_925 ();
 sg13g2_decap_8 FILLER_5_932 ();
 sg13g2_decap_8 FILLER_5_939 ();
 sg13g2_decap_8 FILLER_5_946 ();
 sg13g2_decap_8 FILLER_5_953 ();
 sg13g2_decap_8 FILLER_5_960 ();
 sg13g2_decap_8 FILLER_5_967 ();
 sg13g2_decap_8 FILLER_5_974 ();
 sg13g2_decap_8 FILLER_5_981 ();
 sg13g2_decap_8 FILLER_5_988 ();
 sg13g2_decap_8 FILLER_5_995 ();
 sg13g2_decap_8 FILLER_5_1002 ();
 sg13g2_decap_8 FILLER_5_1009 ();
 sg13g2_decap_8 FILLER_5_1016 ();
 sg13g2_decap_4 FILLER_5_1023 ();
 sg13g2_fill_2 FILLER_5_1027 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_fill_1 FILLER_6_26 ();
 sg13g2_decap_4 FILLER_6_45 ();
 sg13g2_decap_4 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_81 ();
 sg13g2_fill_2 FILLER_6_104 ();
 sg13g2_decap_4 FILLER_6_206 ();
 sg13g2_fill_2 FILLER_6_219 ();
 sg13g2_fill_1 FILLER_6_265 ();
 sg13g2_fill_2 FILLER_6_289 ();
 sg13g2_fill_1 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_351 ();
 sg13g2_fill_2 FILLER_6_361 ();
 sg13g2_fill_2 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_409 ();
 sg13g2_decap_8 FILLER_6_416 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_8 FILLER_6_430 ();
 sg13g2_fill_1 FILLER_6_461 ();
 sg13g2_decap_8 FILLER_6_471 ();
 sg13g2_fill_2 FILLER_6_478 ();
 sg13g2_fill_2 FILLER_6_544 ();
 sg13g2_decap_8 FILLER_6_573 ();
 sg13g2_fill_1 FILLER_6_580 ();
 sg13g2_decap_4 FILLER_6_608 ();
 sg13g2_fill_1 FILLER_6_612 ();
 sg13g2_decap_8 FILLER_6_622 ();
 sg13g2_decap_8 FILLER_6_629 ();
 sg13g2_decap_8 FILLER_6_709 ();
 sg13g2_decap_8 FILLER_6_716 ();
 sg13g2_decap_8 FILLER_6_723 ();
 sg13g2_decap_8 FILLER_6_730 ();
 sg13g2_decap_8 FILLER_6_737 ();
 sg13g2_decap_8 FILLER_6_744 ();
 sg13g2_decap_8 FILLER_6_751 ();
 sg13g2_decap_8 FILLER_6_758 ();
 sg13g2_decap_8 FILLER_6_765 ();
 sg13g2_decap_8 FILLER_6_772 ();
 sg13g2_decap_8 FILLER_6_779 ();
 sg13g2_decap_8 FILLER_6_786 ();
 sg13g2_decap_8 FILLER_6_793 ();
 sg13g2_decap_8 FILLER_6_800 ();
 sg13g2_decap_8 FILLER_6_807 ();
 sg13g2_decap_8 FILLER_6_814 ();
 sg13g2_decap_8 FILLER_6_821 ();
 sg13g2_decap_8 FILLER_6_828 ();
 sg13g2_decap_8 FILLER_6_835 ();
 sg13g2_decap_8 FILLER_6_842 ();
 sg13g2_decap_8 FILLER_6_849 ();
 sg13g2_decap_8 FILLER_6_856 ();
 sg13g2_decap_8 FILLER_6_863 ();
 sg13g2_decap_8 FILLER_6_870 ();
 sg13g2_decap_8 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_6_884 ();
 sg13g2_decap_8 FILLER_6_891 ();
 sg13g2_decap_8 FILLER_6_898 ();
 sg13g2_decap_8 FILLER_6_905 ();
 sg13g2_decap_8 FILLER_6_912 ();
 sg13g2_decap_8 FILLER_6_919 ();
 sg13g2_decap_8 FILLER_6_926 ();
 sg13g2_decap_8 FILLER_6_933 ();
 sg13g2_decap_8 FILLER_6_940 ();
 sg13g2_decap_8 FILLER_6_947 ();
 sg13g2_decap_8 FILLER_6_954 ();
 sg13g2_decap_8 FILLER_6_961 ();
 sg13g2_decap_8 FILLER_6_968 ();
 sg13g2_decap_8 FILLER_6_975 ();
 sg13g2_decap_8 FILLER_6_982 ();
 sg13g2_decap_8 FILLER_6_989 ();
 sg13g2_decap_8 FILLER_6_996 ();
 sg13g2_decap_8 FILLER_6_1003 ();
 sg13g2_decap_8 FILLER_6_1010 ();
 sg13g2_decap_8 FILLER_6_1017 ();
 sg13g2_decap_4 FILLER_6_1024 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_2 ();
 sg13g2_decap_4 FILLER_7_30 ();
 sg13g2_fill_2 FILLER_7_61 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_fill_1 FILLER_7_73 ();
 sg13g2_fill_2 FILLER_7_84 ();
 sg13g2_fill_1 FILLER_7_86 ();
 sg13g2_decap_8 FILLER_7_102 ();
 sg13g2_decap_8 FILLER_7_109 ();
 sg13g2_decap_4 FILLER_7_125 ();
 sg13g2_fill_1 FILLER_7_129 ();
 sg13g2_fill_1 FILLER_7_139 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_decap_4 FILLER_7_193 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_227 ();
 sg13g2_fill_2 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_267 ();
 sg13g2_decap_8 FILLER_7_274 ();
 sg13g2_decap_4 FILLER_7_294 ();
 sg13g2_decap_4 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_fill_2 FILLER_7_372 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_fill_1 FILLER_7_441 ();
 sg13g2_fill_2 FILLER_7_495 ();
 sg13g2_decap_8 FILLER_7_510 ();
 sg13g2_fill_1 FILLER_7_521 ();
 sg13g2_fill_1 FILLER_7_530 ();
 sg13g2_decap_8 FILLER_7_545 ();
 sg13g2_decap_8 FILLER_7_552 ();
 sg13g2_fill_2 FILLER_7_581 ();
 sg13g2_fill_1 FILLER_7_583 ();
 sg13g2_fill_1 FILLER_7_593 ();
 sg13g2_decap_4 FILLER_7_598 ();
 sg13g2_fill_2 FILLER_7_611 ();
 sg13g2_fill_1 FILLER_7_613 ();
 sg13g2_decap_4 FILLER_7_673 ();
 sg13g2_fill_2 FILLER_7_687 ();
 sg13g2_fill_1 FILLER_7_689 ();
 sg13g2_decap_8 FILLER_7_712 ();
 sg13g2_decap_8 FILLER_7_719 ();
 sg13g2_decap_8 FILLER_7_726 ();
 sg13g2_decap_8 FILLER_7_733 ();
 sg13g2_decap_8 FILLER_7_740 ();
 sg13g2_decap_8 FILLER_7_747 ();
 sg13g2_decap_8 FILLER_7_754 ();
 sg13g2_decap_8 FILLER_7_761 ();
 sg13g2_decap_8 FILLER_7_768 ();
 sg13g2_decap_8 FILLER_7_775 ();
 sg13g2_decap_8 FILLER_7_782 ();
 sg13g2_decap_8 FILLER_7_789 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_decap_8 FILLER_7_803 ();
 sg13g2_decap_8 FILLER_7_810 ();
 sg13g2_decap_8 FILLER_7_817 ();
 sg13g2_decap_8 FILLER_7_824 ();
 sg13g2_decap_4 FILLER_7_831 ();
 sg13g2_fill_1 FILLER_7_839 ();
 sg13g2_decap_8 FILLER_7_850 ();
 sg13g2_decap_8 FILLER_7_857 ();
 sg13g2_decap_8 FILLER_7_864 ();
 sg13g2_decap_8 FILLER_7_871 ();
 sg13g2_decap_8 FILLER_7_878 ();
 sg13g2_decap_8 FILLER_7_885 ();
 sg13g2_decap_8 FILLER_7_892 ();
 sg13g2_decap_8 FILLER_7_899 ();
 sg13g2_decap_8 FILLER_7_906 ();
 sg13g2_decap_8 FILLER_7_913 ();
 sg13g2_decap_8 FILLER_7_920 ();
 sg13g2_decap_8 FILLER_7_927 ();
 sg13g2_decap_8 FILLER_7_934 ();
 sg13g2_decap_8 FILLER_7_941 ();
 sg13g2_decap_8 FILLER_7_948 ();
 sg13g2_decap_8 FILLER_7_955 ();
 sg13g2_decap_8 FILLER_7_962 ();
 sg13g2_decap_8 FILLER_7_969 ();
 sg13g2_decap_8 FILLER_7_976 ();
 sg13g2_decap_8 FILLER_7_983 ();
 sg13g2_decap_8 FILLER_7_990 ();
 sg13g2_decap_8 FILLER_7_997 ();
 sg13g2_decap_8 FILLER_7_1004 ();
 sg13g2_decap_8 FILLER_7_1011 ();
 sg13g2_decap_8 FILLER_7_1018 ();
 sg13g2_decap_4 FILLER_7_1025 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_30 ();
 sg13g2_fill_2 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_58 ();
 sg13g2_fill_2 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_163 ();
 sg13g2_fill_2 FILLER_8_177 ();
 sg13g2_fill_1 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_fill_2 FILLER_8_248 ();
 sg13g2_fill_1 FILLER_8_250 ();
 sg13g2_decap_8 FILLER_8_269 ();
 sg13g2_decap_8 FILLER_8_276 ();
 sg13g2_fill_2 FILLER_8_283 ();
 sg13g2_fill_1 FILLER_8_285 ();
 sg13g2_fill_1 FILLER_8_291 ();
 sg13g2_fill_2 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_339 ();
 sg13g2_decap_8 FILLER_8_346 ();
 sg13g2_fill_2 FILLER_8_380 ();
 sg13g2_fill_1 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_fill_1 FILLER_8_430 ();
 sg13g2_fill_1 FILLER_8_452 ();
 sg13g2_fill_1 FILLER_8_468 ();
 sg13g2_decap_8 FILLER_8_479 ();
 sg13g2_decap_8 FILLER_8_486 ();
 sg13g2_decap_4 FILLER_8_493 ();
 sg13g2_fill_2 FILLER_8_524 ();
 sg13g2_fill_2 FILLER_8_531 ();
 sg13g2_fill_1 FILLER_8_533 ();
 sg13g2_decap_4 FILLER_8_548 ();
 sg13g2_fill_1 FILLER_8_552 ();
 sg13g2_fill_1 FILLER_8_653 ();
 sg13g2_decap_8 FILLER_8_681 ();
 sg13g2_fill_1 FILLER_8_688 ();
 sg13g2_decap_8 FILLER_8_717 ();
 sg13g2_decap_8 FILLER_8_724 ();
 sg13g2_decap_8 FILLER_8_731 ();
 sg13g2_decap_4 FILLER_8_738 ();
 sg13g2_fill_1 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_748 ();
 sg13g2_decap_8 FILLER_8_755 ();
 sg13g2_decap_8 FILLER_8_762 ();
 sg13g2_decap_8 FILLER_8_769 ();
 sg13g2_decap_8 FILLER_8_776 ();
 sg13g2_decap_8 FILLER_8_783 ();
 sg13g2_decap_4 FILLER_8_790 ();
 sg13g2_fill_1 FILLER_8_802 ();
 sg13g2_decap_4 FILLER_8_822 ();
 sg13g2_fill_2 FILLER_8_826 ();
 sg13g2_fill_2 FILLER_8_842 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_decap_8 FILLER_8_875 ();
 sg13g2_decap_8 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_889 ();
 sg13g2_decap_8 FILLER_8_896 ();
 sg13g2_decap_8 FILLER_8_903 ();
 sg13g2_decap_8 FILLER_8_910 ();
 sg13g2_decap_8 FILLER_8_917 ();
 sg13g2_decap_8 FILLER_8_924 ();
 sg13g2_decap_8 FILLER_8_931 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_945 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_8 FILLER_8_959 ();
 sg13g2_decap_8 FILLER_8_966 ();
 sg13g2_decap_8 FILLER_8_973 ();
 sg13g2_decap_8 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_decap_8 FILLER_8_994 ();
 sg13g2_decap_8 FILLER_8_1001 ();
 sg13g2_decap_8 FILLER_8_1008 ();
 sg13g2_decap_8 FILLER_8_1015 ();
 sg13g2_decap_8 FILLER_8_1022 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_1 FILLER_9_39 ();
 sg13g2_fill_1 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_63 ();
 sg13g2_fill_1 FILLER_9_65 ();
 sg13g2_fill_2 FILLER_9_75 ();
 sg13g2_fill_1 FILLER_9_77 ();
 sg13g2_fill_1 FILLER_9_167 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_268 ();
 sg13g2_decap_4 FILLER_9_279 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_355 ();
 sg13g2_fill_2 FILLER_9_397 ();
 sg13g2_fill_2 FILLER_9_408 ();
 sg13g2_decap_4 FILLER_9_454 ();
 sg13g2_decap_8 FILLER_9_478 ();
 sg13g2_fill_2 FILLER_9_485 ();
 sg13g2_decap_8 FILLER_9_491 ();
 sg13g2_decap_4 FILLER_9_498 ();
 sg13g2_fill_1 FILLER_9_502 ();
 sg13g2_decap_8 FILLER_9_509 ();
 sg13g2_decap_8 FILLER_9_516 ();
 sg13g2_decap_4 FILLER_9_523 ();
 sg13g2_fill_1 FILLER_9_527 ();
 sg13g2_fill_2 FILLER_9_548 ();
 sg13g2_fill_2 FILLER_9_560 ();
 sg13g2_decap_4 FILLER_9_576 ();
 sg13g2_decap_8 FILLER_9_593 ();
 sg13g2_fill_1 FILLER_9_600 ();
 sg13g2_decap_4 FILLER_9_609 ();
 sg13g2_fill_1 FILLER_9_627 ();
 sg13g2_fill_1 FILLER_9_643 ();
 sg13g2_fill_1 FILLER_9_648 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_fill_2 FILLER_9_665 ();
 sg13g2_decap_4 FILLER_9_714 ();
 sg13g2_fill_2 FILLER_9_718 ();
 sg13g2_decap_4 FILLER_9_733 ();
 sg13g2_decap_4 FILLER_9_765 ();
 sg13g2_fill_1 FILLER_9_769 ();
 sg13g2_fill_1 FILLER_9_829 ();
 sg13g2_decap_8 FILLER_9_866 ();
 sg13g2_decap_8 FILLER_9_873 ();
 sg13g2_fill_2 FILLER_9_880 ();
 sg13g2_decap_8 FILLER_9_885 ();
 sg13g2_fill_2 FILLER_9_892 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_fill_2 FILLER_10_31 ();
 sg13g2_fill_1 FILLER_10_33 ();
 sg13g2_decap_8 FILLER_10_125 ();
 sg13g2_decap_4 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_149 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_decap_4 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_fill_1 FILLER_10_221 ();
 sg13g2_fill_2 FILLER_10_245 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_fill_2 FILLER_10_297 ();
 sg13g2_fill_1 FILLER_10_326 ();
 sg13g2_decap_4 FILLER_10_336 ();
 sg13g2_fill_1 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_fill_2 FILLER_10_386 ();
 sg13g2_fill_2 FILLER_10_417 ();
 sg13g2_fill_1 FILLER_10_419 ();
 sg13g2_fill_2 FILLER_10_435 ();
 sg13g2_fill_1 FILLER_10_437 ();
 sg13g2_fill_1 FILLER_10_446 ();
 sg13g2_fill_2 FILLER_10_452 ();
 sg13g2_fill_2 FILLER_10_476 ();
 sg13g2_fill_2 FILLER_10_484 ();
 sg13g2_fill_1 FILLER_10_486 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_fill_2 FILLER_10_525 ();
 sg13g2_fill_1 FILLER_10_527 ();
 sg13g2_decap_4 FILLER_10_532 ();
 sg13g2_fill_1 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_540 ();
 sg13g2_decap_8 FILLER_10_547 ();
 sg13g2_fill_2 FILLER_10_554 ();
 sg13g2_fill_1 FILLER_10_556 ();
 sg13g2_fill_2 FILLER_10_588 ();
 sg13g2_fill_2 FILLER_10_612 ();
 sg13g2_fill_1 FILLER_10_614 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_4 FILLER_10_651 ();
 sg13g2_fill_1 FILLER_10_682 ();
 sg13g2_decap_4 FILLER_10_706 ();
 sg13g2_fill_2 FILLER_10_738 ();
 sg13g2_fill_1 FILLER_10_740 ();
 sg13g2_decap_8 FILLER_10_783 ();
 sg13g2_fill_1 FILLER_10_790 ();
 sg13g2_fill_2 FILLER_10_796 ();
 sg13g2_fill_1 FILLER_10_835 ();
 sg13g2_fill_1 FILLER_10_876 ();
 sg13g2_decap_8 FILLER_10_904 ();
 sg13g2_decap_8 FILLER_10_911 ();
 sg13g2_decap_8 FILLER_10_918 ();
 sg13g2_decap_8 FILLER_10_925 ();
 sg13g2_decap_8 FILLER_10_932 ();
 sg13g2_decap_8 FILLER_10_939 ();
 sg13g2_decap_8 FILLER_10_946 ();
 sg13g2_decap_8 FILLER_10_953 ();
 sg13g2_decap_8 FILLER_10_960 ();
 sg13g2_decap_8 FILLER_10_967 ();
 sg13g2_decap_8 FILLER_10_974 ();
 sg13g2_decap_8 FILLER_10_981 ();
 sg13g2_decap_8 FILLER_10_988 ();
 sg13g2_decap_8 FILLER_10_995 ();
 sg13g2_decap_8 FILLER_10_1002 ();
 sg13g2_decap_8 FILLER_10_1009 ();
 sg13g2_decap_8 FILLER_10_1016 ();
 sg13g2_decap_4 FILLER_10_1023 ();
 sg13g2_fill_2 FILLER_10_1027 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_58 ();
 sg13g2_decap_4 FILLER_11_65 ();
 sg13g2_fill_1 FILLER_11_74 ();
 sg13g2_decap_4 FILLER_11_114 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_decap_8 FILLER_11_136 ();
 sg13g2_decap_8 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_decap_4 FILLER_11_212 ();
 sg13g2_decap_4 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_8 FILLER_11_320 ();
 sg13g2_fill_2 FILLER_11_327 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_fill_2 FILLER_11_362 ();
 sg13g2_fill_1 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_411 ();
 sg13g2_fill_2 FILLER_11_418 ();
 sg13g2_fill_1 FILLER_11_420 ();
 sg13g2_fill_1 FILLER_11_436 ();
 sg13g2_fill_1 FILLER_11_443 ();
 sg13g2_decap_8 FILLER_11_450 ();
 sg13g2_decap_4 FILLER_11_457 ();
 sg13g2_fill_1 FILLER_11_461 ();
 sg13g2_decap_4 FILLER_11_476 ();
 sg13g2_fill_1 FILLER_11_480 ();
 sg13g2_fill_2 FILLER_11_491 ();
 sg13g2_fill_1 FILLER_11_493 ();
 sg13g2_fill_1 FILLER_11_499 ();
 sg13g2_decap_8 FILLER_11_509 ();
 sg13g2_decap_4 FILLER_11_516 ();
 sg13g2_fill_1 FILLER_11_520 ();
 sg13g2_decap_4 FILLER_11_552 ();
 sg13g2_fill_2 FILLER_11_576 ();
 sg13g2_fill_1 FILLER_11_578 ();
 sg13g2_fill_2 FILLER_11_651 ();
 sg13g2_fill_1 FILLER_11_653 ();
 sg13g2_fill_2 FILLER_11_689 ();
 sg13g2_fill_1 FILLER_11_691 ();
 sg13g2_decap_8 FILLER_11_701 ();
 sg13g2_decap_4 FILLER_11_708 ();
 sg13g2_fill_1 FILLER_11_769 ();
 sg13g2_fill_2 FILLER_11_792 ();
 sg13g2_fill_1 FILLER_11_794 ();
 sg13g2_fill_2 FILLER_11_808 ();
 sg13g2_fill_2 FILLER_11_821 ();
 sg13g2_fill_2 FILLER_11_832 ();
 sg13g2_fill_2 FILLER_11_839 ();
 sg13g2_fill_1 FILLER_11_881 ();
 sg13g2_decap_8 FILLER_11_917 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_decap_8 FILLER_11_945 ();
 sg13g2_decap_8 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_8 FILLER_11_1001 ();
 sg13g2_decap_8 FILLER_11_1008 ();
 sg13g2_decap_8 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1022 ();
 sg13g2_decap_4 FILLER_12_59 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_83 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_108 ();
 sg13g2_fill_2 FILLER_12_149 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_fill_2 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_219 ();
 sg13g2_decap_4 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_decap_4 FILLER_12_291 ();
 sg13g2_fill_2 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_324 ();
 sg13g2_fill_2 FILLER_12_375 ();
 sg13g2_fill_1 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_fill_1 FILLER_12_417 ();
 sg13g2_decap_8 FILLER_12_449 ();
 sg13g2_decap_4 FILLER_12_456 ();
 sg13g2_fill_1 FILLER_12_460 ();
 sg13g2_fill_2 FILLER_12_485 ();
 sg13g2_fill_2 FILLER_12_510 ();
 sg13g2_decap_4 FILLER_12_540 ();
 sg13g2_fill_1 FILLER_12_544 ();
 sg13g2_decap_4 FILLER_12_558 ();
 sg13g2_fill_2 FILLER_12_589 ();
 sg13g2_fill_1 FILLER_12_591 ();
 sg13g2_decap_4 FILLER_12_609 ();
 sg13g2_decap_4 FILLER_12_622 ();
 sg13g2_decap_8 FILLER_12_642 ();
 sg13g2_fill_2 FILLER_12_649 ();
 sg13g2_fill_1 FILLER_12_651 ();
 sg13g2_fill_2 FILLER_12_669 ();
 sg13g2_fill_1 FILLER_12_671 ();
 sg13g2_fill_2 FILLER_12_748 ();
 sg13g2_fill_2 FILLER_12_754 ();
 sg13g2_fill_2 FILLER_12_783 ();
 sg13g2_fill_2 FILLER_12_793 ();
 sg13g2_fill_2 FILLER_12_827 ();
 sg13g2_fill_1 FILLER_12_829 ();
 sg13g2_fill_2 FILLER_12_848 ();
 sg13g2_fill_1 FILLER_12_850 ();
 sg13g2_decap_8 FILLER_12_878 ();
 sg13g2_fill_2 FILLER_12_885 ();
 sg13g2_fill_1 FILLER_12_887 ();
 sg13g2_decap_8 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_909 ();
 sg13g2_decap_8 FILLER_12_916 ();
 sg13g2_decap_8 FILLER_12_923 ();
 sg13g2_decap_8 FILLER_12_930 ();
 sg13g2_decap_8 FILLER_12_937 ();
 sg13g2_decap_8 FILLER_12_944 ();
 sg13g2_decap_8 FILLER_12_951 ();
 sg13g2_decap_8 FILLER_12_958 ();
 sg13g2_decap_8 FILLER_12_965 ();
 sg13g2_decap_8 FILLER_12_972 ();
 sg13g2_decap_8 FILLER_12_979 ();
 sg13g2_decap_8 FILLER_12_986 ();
 sg13g2_decap_8 FILLER_12_993 ();
 sg13g2_decap_8 FILLER_12_1000 ();
 sg13g2_decap_8 FILLER_12_1007 ();
 sg13g2_decap_8 FILLER_12_1014 ();
 sg13g2_decap_4 FILLER_12_1021 ();
 sg13g2_fill_1 FILLER_13_8 ();
 sg13g2_fill_2 FILLER_13_22 ();
 sg13g2_fill_1 FILLER_13_24 ();
 sg13g2_fill_2 FILLER_13_38 ();
 sg13g2_decap_8 FILLER_13_54 ();
 sg13g2_fill_1 FILLER_13_61 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_118 ();
 sg13g2_fill_1 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_174 ();
 sg13g2_fill_2 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_187 ();
 sg13g2_fill_1 FILLER_13_189 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_223 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_decap_4 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_241 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_254 ();
 sg13g2_decap_8 FILLER_13_328 ();
 sg13g2_fill_2 FILLER_13_335 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_4 FILLER_13_354 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_13_409 ();
 sg13g2_fill_1 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_4 FILLER_13_448 ();
 sg13g2_fill_1 FILLER_13_452 ();
 sg13g2_fill_2 FILLER_13_477 ();
 sg13g2_fill_2 FILLER_13_487 ();
 sg13g2_decap_8 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_537 ();
 sg13g2_decap_8 FILLER_13_544 ();
 sg13g2_decap_4 FILLER_13_564 ();
 sg13g2_decap_8 FILLER_13_573 ();
 sg13g2_decap_8 FILLER_13_580 ();
 sg13g2_decap_8 FILLER_13_587 ();
 sg13g2_decap_8 FILLER_13_597 ();
 sg13g2_decap_8 FILLER_13_604 ();
 sg13g2_decap_8 FILLER_13_611 ();
 sg13g2_decap_4 FILLER_13_618 ();
 sg13g2_fill_1 FILLER_13_635 ();
 sg13g2_fill_1 FILLER_13_662 ();
 sg13g2_fill_2 FILLER_13_668 ();
 sg13g2_fill_1 FILLER_13_670 ();
 sg13g2_fill_2 FILLER_13_684 ();
 sg13g2_decap_8 FILLER_13_694 ();
 sg13g2_decap_8 FILLER_13_701 ();
 sg13g2_decap_8 FILLER_13_708 ();
 sg13g2_decap_8 FILLER_13_715 ();
 sg13g2_fill_2 FILLER_13_722 ();
 sg13g2_fill_2 FILLER_13_748 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_4 FILLER_13_770 ();
 sg13g2_fill_1 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_fill_1 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_827 ();
 sg13g2_fill_2 FILLER_13_834 ();
 sg13g2_fill_1 FILLER_13_836 ();
 sg13g2_decap_8 FILLER_13_915 ();
 sg13g2_decap_8 FILLER_13_922 ();
 sg13g2_decap_8 FILLER_13_929 ();
 sg13g2_decap_8 FILLER_13_936 ();
 sg13g2_decap_8 FILLER_13_943 ();
 sg13g2_decap_8 FILLER_13_950 ();
 sg13g2_decap_8 FILLER_13_957 ();
 sg13g2_decap_8 FILLER_13_964 ();
 sg13g2_decap_8 FILLER_13_971 ();
 sg13g2_decap_8 FILLER_13_978 ();
 sg13g2_decap_8 FILLER_13_985 ();
 sg13g2_decap_8 FILLER_13_992 ();
 sg13g2_decap_8 FILLER_13_999 ();
 sg13g2_decap_8 FILLER_13_1006 ();
 sg13g2_decap_8 FILLER_13_1013 ();
 sg13g2_decap_8 FILLER_13_1020 ();
 sg13g2_fill_2 FILLER_13_1027 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_decap_4 FILLER_14_81 ();
 sg13g2_fill_2 FILLER_14_85 ();
 sg13g2_fill_2 FILLER_14_100 ();
 sg13g2_fill_1 FILLER_14_117 ();
 sg13g2_decap_4 FILLER_14_127 ();
 sg13g2_decap_8 FILLER_14_135 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_188 ();
 sg13g2_decap_4 FILLER_14_221 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_4 FILLER_14_257 ();
 sg13g2_fill_2 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_fill_2 FILLER_14_323 ();
 sg13g2_fill_1 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_367 ();
 sg13g2_decap_4 FILLER_14_374 ();
 sg13g2_fill_2 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_fill_1 FILLER_14_418 ();
 sg13g2_fill_1 FILLER_14_443 ();
 sg13g2_decap_8 FILLER_14_450 ();
 sg13g2_decap_4 FILLER_14_470 ();
 sg13g2_decap_8 FILLER_14_501 ();
 sg13g2_decap_8 FILLER_14_508 ();
 sg13g2_fill_2 FILLER_14_515 ();
 sg13g2_fill_1 FILLER_14_517 ();
 sg13g2_decap_8 FILLER_14_530 ();
 sg13g2_decap_4 FILLER_14_537 ();
 sg13g2_fill_2 FILLER_14_541 ();
 sg13g2_decap_8 FILLER_14_549 ();
 sg13g2_fill_1 FILLER_14_556 ();
 sg13g2_fill_2 FILLER_14_570 ();
 sg13g2_decap_4 FILLER_14_586 ();
 sg13g2_fill_1 FILLER_14_632 ();
 sg13g2_fill_1 FILLER_14_641 ();
 sg13g2_decap_8 FILLER_14_710 ();
 sg13g2_decap_4 FILLER_14_717 ();
 sg13g2_fill_1 FILLER_14_721 ();
 sg13g2_fill_2 FILLER_14_752 ();
 sg13g2_fill_1 FILLER_14_754 ();
 sg13g2_decap_4 FILLER_14_769 ();
 sg13g2_decap_4 FILLER_14_790 ();
 sg13g2_fill_1 FILLER_14_794 ();
 sg13g2_decap_4 FILLER_14_827 ();
 sg13g2_fill_1 FILLER_14_831 ();
 sg13g2_decap_4 FILLER_14_873 ();
 sg13g2_fill_2 FILLER_14_877 ();
 sg13g2_decap_8 FILLER_14_882 ();
 sg13g2_decap_8 FILLER_14_889 ();
 sg13g2_fill_1 FILLER_14_896 ();
 sg13g2_decap_8 FILLER_14_960 ();
 sg13g2_fill_2 FILLER_14_967 ();
 sg13g2_fill_1 FILLER_14_969 ();
 sg13g2_decap_4 FILLER_14_974 ();
 sg13g2_fill_1 FILLER_14_978 ();
 sg13g2_decap_8 FILLER_14_988 ();
 sg13g2_decap_8 FILLER_14_995 ();
 sg13g2_decap_8 FILLER_14_1002 ();
 sg13g2_decap_8 FILLER_14_1009 ();
 sg13g2_decap_8 FILLER_14_1016 ();
 sg13g2_decap_4 FILLER_14_1023 ();
 sg13g2_fill_2 FILLER_14_1027 ();
 sg13g2_decap_4 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_8 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_fill_2 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_79 ();
 sg13g2_fill_2 FILLER_15_86 ();
 sg13g2_fill_2 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_117 ();
 sg13g2_fill_2 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_156 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_213 ();
 sg13g2_decap_4 FILLER_15_222 ();
 sg13g2_decap_4 FILLER_15_262 ();
 sg13g2_fill_2 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_1 FILLER_15_338 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_fill_2 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_15_414 ();
 sg13g2_fill_1 FILLER_15_416 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_2 FILLER_15_458 ();
 sg13g2_decap_8 FILLER_15_465 ();
 sg13g2_fill_2 FILLER_15_472 ();
 sg13g2_fill_1 FILLER_15_474 ();
 sg13g2_fill_1 FILLER_15_495 ();
 sg13g2_decap_4 FILLER_15_505 ();
 sg13g2_fill_2 FILLER_15_518 ();
 sg13g2_fill_1 FILLER_15_520 ();
 sg13g2_fill_1 FILLER_15_531 ();
 sg13g2_fill_1 FILLER_15_559 ();
 sg13g2_fill_2 FILLER_15_587 ();
 sg13g2_decap_8 FILLER_15_617 ();
 sg13g2_fill_1 FILLER_15_624 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_4 FILLER_15_665 ();
 sg13g2_decap_4 FILLER_15_687 ();
 sg13g2_fill_2 FILLER_15_691 ();
 sg13g2_fill_2 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_820 ();
 sg13g2_fill_1 FILLER_15_827 ();
 sg13g2_fill_2 FILLER_15_849 ();
 sg13g2_fill_1 FILLER_15_851 ();
 sg13g2_decap_4 FILLER_15_902 ();
 sg13g2_fill_1 FILLER_15_906 ();
 sg13g2_decap_8 FILLER_15_920 ();
 sg13g2_decap_8 FILLER_15_927 ();
 sg13g2_fill_2 FILLER_15_934 ();
 sg13g2_decap_8 FILLER_15_998 ();
 sg13g2_decap_8 FILLER_15_1005 ();
 sg13g2_decap_8 FILLER_15_1012 ();
 sg13g2_decap_8 FILLER_15_1019 ();
 sg13g2_fill_2 FILLER_15_1026 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_4 FILLER_16_11 ();
 sg13g2_fill_1 FILLER_16_33 ();
 sg13g2_fill_2 FILLER_16_40 ();
 sg13g2_fill_1 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_48 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_decap_4 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_decap_8 FILLER_16_260 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_4 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_348 ();
 sg13g2_fill_2 FILLER_16_359 ();
 sg13g2_decap_4 FILLER_16_376 ();
 sg13g2_fill_2 FILLER_16_380 ();
 sg13g2_fill_1 FILLER_16_391 ();
 sg13g2_fill_1 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_4 FILLER_16_419 ();
 sg13g2_fill_2 FILLER_16_423 ();
 sg13g2_decap_8 FILLER_16_435 ();
 sg13g2_decap_8 FILLER_16_442 ();
 sg13g2_decap_8 FILLER_16_468 ();
 sg13g2_decap_4 FILLER_16_475 ();
 sg13g2_decap_8 FILLER_16_545 ();
 sg13g2_fill_1 FILLER_16_552 ();
 sg13g2_fill_2 FILLER_16_576 ();
 sg13g2_fill_1 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_599 ();
 sg13g2_fill_2 FILLER_16_606 ();
 sg13g2_fill_2 FILLER_16_638 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_fill_2 FILLER_16_707 ();
 sg13g2_fill_1 FILLER_16_709 ();
 sg13g2_fill_2 FILLER_16_715 ();
 sg13g2_fill_1 FILLER_16_761 ();
 sg13g2_decap_4 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_fill_2 FILLER_16_833 ();
 sg13g2_fill_1 FILLER_16_835 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_decap_8 FILLER_16_875 ();
 sg13g2_fill_2 FILLER_16_882 ();
 sg13g2_fill_1 FILLER_16_884 ();
 sg13g2_fill_2 FILLER_16_917 ();
 sg13g2_fill_1 FILLER_16_969 ();
 sg13g2_decap_8 FILLER_16_1002 ();
 sg13g2_decap_8 FILLER_16_1009 ();
 sg13g2_decap_8 FILLER_16_1016 ();
 sg13g2_decap_4 FILLER_16_1023 ();
 sg13g2_fill_2 FILLER_16_1027 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_6 ();
 sg13g2_decap_4 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_90 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_1 FILLER_17_204 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_fill_1 FILLER_17_338 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_fill_2 FILLER_17_383 ();
 sg13g2_fill_1 FILLER_17_385 ();
 sg13g2_decap_4 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_395 ();
 sg13g2_decap_4 FILLER_17_413 ();
 sg13g2_fill_2 FILLER_17_423 ();
 sg13g2_fill_1 FILLER_17_425 ();
 sg13g2_decap_8 FILLER_17_444 ();
 sg13g2_fill_1 FILLER_17_451 ();
 sg13g2_fill_1 FILLER_17_457 ();
 sg13g2_decap_8 FILLER_17_463 ();
 sg13g2_decap_4 FILLER_17_470 ();
 sg13g2_decap_4 FILLER_17_478 ();
 sg13g2_decap_8 FILLER_17_492 ();
 sg13g2_decap_8 FILLER_17_499 ();
 sg13g2_decap_8 FILLER_17_506 ();
 sg13g2_decap_4 FILLER_17_513 ();
 sg13g2_fill_1 FILLER_17_517 ();
 sg13g2_decap_4 FILLER_17_528 ();
 sg13g2_fill_1 FILLER_17_541 ();
 sg13g2_decap_8 FILLER_17_551 ();
 sg13g2_decap_4 FILLER_17_558 ();
 sg13g2_fill_1 FILLER_17_562 ();
 sg13g2_fill_2 FILLER_17_600 ();
 sg13g2_decap_8 FILLER_17_618 ();
 sg13g2_fill_2 FILLER_17_625 ();
 sg13g2_fill_1 FILLER_17_627 ();
 sg13g2_fill_2 FILLER_17_676 ();
 sg13g2_fill_1 FILLER_17_678 ();
 sg13g2_decap_4 FILLER_17_719 ();
 sg13g2_fill_1 FILLER_17_788 ();
 sg13g2_fill_2 FILLER_17_807 ();
 sg13g2_fill_2 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_838 ();
 sg13g2_fill_1 FILLER_17_845 ();
 sg13g2_fill_2 FILLER_17_855 ();
 sg13g2_fill_1 FILLER_17_857 ();
 sg13g2_decap_8 FILLER_17_871 ();
 sg13g2_fill_1 FILLER_17_878 ();
 sg13g2_fill_1 FILLER_17_901 ();
 sg13g2_fill_2 FILLER_17_972 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_fill_2 FILLER_18_4 ();
 sg13g2_fill_1 FILLER_18_6 ();
 sg13g2_fill_2 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_80 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_decap_4 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_fill_2 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_251 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_decap_4 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_321 ();
 sg13g2_fill_2 FILLER_18_332 ();
 sg13g2_decap_4 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_decap_4 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_414 ();
 sg13g2_decap_4 FILLER_18_444 ();
 sg13g2_fill_1 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_459 ();
 sg13g2_fill_1 FILLER_18_478 ();
 sg13g2_decap_8 FILLER_18_496 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_fill_2 FILLER_18_567 ();
 sg13g2_fill_1 FILLER_18_569 ();
 sg13g2_decap_8 FILLER_18_585 ();
 sg13g2_fill_2 FILLER_18_592 ();
 sg13g2_fill_2 FILLER_18_599 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_fill_1 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_646 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_4 FILLER_18_665 ();
 sg13g2_fill_1 FILLER_18_669 ();
 sg13g2_fill_2 FILLER_18_675 ();
 sg13g2_fill_2 FILLER_18_690 ();
 sg13g2_fill_1 FILLER_18_692 ();
 sg13g2_decap_4 FILLER_18_702 ();
 sg13g2_fill_1 FILLER_18_706 ();
 sg13g2_decap_4 FILLER_18_720 ();
 sg13g2_fill_2 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_fill_2 FILLER_18_810 ();
 sg13g2_decap_8 FILLER_18_846 ();
 sg13g2_fill_1 FILLER_18_853 ();
 sg13g2_fill_1 FILLER_18_894 ();
 sg13g2_fill_1 FILLER_18_904 ();
 sg13g2_fill_2 FILLER_18_919 ();
 sg13g2_decap_8 FILLER_18_930 ();
 sg13g2_decap_8 FILLER_18_937 ();
 sg13g2_fill_2 FILLER_18_944 ();
 sg13g2_decap_8 FILLER_18_951 ();
 sg13g2_decap_8 FILLER_18_958 ();
 sg13g2_fill_2 FILLER_18_965 ();
 sg13g2_decap_4 FILLER_18_979 ();
 sg13g2_decap_8 FILLER_18_1000 ();
 sg13g2_decap_8 FILLER_18_1007 ();
 sg13g2_decap_8 FILLER_18_1014 ();
 sg13g2_decap_8 FILLER_18_1021 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_fill_1 FILLER_19_52 ();
 sg13g2_decap_4 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_decap_4 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_167 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_1 FILLER_19_258 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_decap_4 FILLER_19_371 ();
 sg13g2_fill_2 FILLER_19_375 ();
 sg13g2_fill_2 FILLER_19_397 ();
 sg13g2_decap_8 FILLER_19_404 ();
 sg13g2_decap_8 FILLER_19_411 ();
 sg13g2_decap_4 FILLER_19_423 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_2 FILLER_19_457 ();
 sg13g2_fill_1 FILLER_19_459 ();
 sg13g2_fill_1 FILLER_19_465 ();
 sg13g2_decap_8 FILLER_19_475 ();
 sg13g2_decap_4 FILLER_19_482 ();
 sg13g2_fill_1 FILLER_19_486 ();
 sg13g2_decap_4 FILLER_19_493 ();
 sg13g2_fill_2 FILLER_19_497 ();
 sg13g2_fill_2 FILLER_19_512 ();
 sg13g2_fill_1 FILLER_19_565 ();
 sg13g2_decap_8 FILLER_19_576 ();
 sg13g2_decap_8 FILLER_19_583 ();
 sg13g2_decap_4 FILLER_19_590 ();
 sg13g2_fill_2 FILLER_19_602 ();
 sg13g2_fill_2 FILLER_19_636 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_fill_1 FILLER_19_663 ();
 sg13g2_fill_2 FILLER_19_674 ();
 sg13g2_fill_1 FILLER_19_676 ();
 sg13g2_fill_2 FILLER_19_690 ();
 sg13g2_fill_1 FILLER_19_739 ();
 sg13g2_fill_2 FILLER_19_757 ();
 sg13g2_fill_1 FILLER_19_759 ();
 sg13g2_decap_4 FILLER_19_769 ();
 sg13g2_fill_1 FILLER_19_773 ();
 sg13g2_fill_2 FILLER_19_841 ();
 sg13g2_fill_1 FILLER_19_843 ();
 sg13g2_fill_2 FILLER_19_851 ();
 sg13g2_fill_2 FILLER_19_866 ();
 sg13g2_decap_8 FILLER_19_877 ();
 sg13g2_decap_8 FILLER_19_884 ();
 sg13g2_fill_2 FILLER_19_917 ();
 sg13g2_fill_1 FILLER_19_919 ();
 sg13g2_fill_1 FILLER_19_929 ();
 sg13g2_decap_8 FILLER_19_957 ();
 sg13g2_decap_8 FILLER_19_964 ();
 sg13g2_fill_2 FILLER_19_971 ();
 sg13g2_decap_8 FILLER_19_1009 ();
 sg13g2_decap_8 FILLER_19_1016 ();
 sg13g2_decap_4 FILLER_19_1023 ();
 sg13g2_fill_2 FILLER_19_1027 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_159 ();
 sg13g2_fill_2 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_241 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_decap_4 FILLER_20_262 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_fill_2 FILLER_20_414 ();
 sg13g2_decap_4 FILLER_20_422 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_fill_1 FILLER_20_441 ();
 sg13g2_fill_1 FILLER_20_472 ();
 sg13g2_decap_8 FILLER_20_478 ();
 sg13g2_fill_2 FILLER_20_485 ();
 sg13g2_fill_1 FILLER_20_487 ();
 sg13g2_fill_2 FILLER_20_501 ();
 sg13g2_fill_1 FILLER_20_503 ();
 sg13g2_decap_4 FILLER_20_541 ();
 sg13g2_fill_2 FILLER_20_554 ();
 sg13g2_fill_1 FILLER_20_556 ();
 sg13g2_decap_8 FILLER_20_597 ();
 sg13g2_fill_2 FILLER_20_604 ();
 sg13g2_decap_8 FILLER_20_610 ();
 sg13g2_decap_8 FILLER_20_617 ();
 sg13g2_fill_2 FILLER_20_624 ();
 sg13g2_fill_1 FILLER_20_626 ();
 sg13g2_fill_2 FILLER_20_637 ();
 sg13g2_fill_2 FILLER_20_655 ();
 sg13g2_fill_1 FILLER_20_657 ();
 sg13g2_fill_2 FILLER_20_712 ();
 sg13g2_fill_1 FILLER_20_733 ();
 sg13g2_decap_8 FILLER_20_761 ();
 sg13g2_decap_8 FILLER_20_768 ();
 sg13g2_fill_1 FILLER_20_775 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_fill_1 FILLER_20_799 ();
 sg13g2_fill_1 FILLER_20_825 ();
 sg13g2_fill_2 FILLER_20_862 ();
 sg13g2_fill_1 FILLER_20_897 ();
 sg13g2_fill_2 FILLER_20_907 ();
 sg13g2_fill_1 FILLER_20_909 ();
 sg13g2_fill_2 FILLER_20_976 ();
 sg13g2_fill_1 FILLER_20_978 ();
 sg13g2_decap_8 FILLER_20_1015 ();
 sg13g2_decap_8 FILLER_20_1022 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_fill_1 FILLER_21_64 ();
 sg13g2_decap_8 FILLER_21_97 ();
 sg13g2_fill_2 FILLER_21_104 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_fill_2 FILLER_21_130 ();
 sg13g2_fill_2 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_143 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_264 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_fill_1 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_4 FILLER_21_417 ();
 sg13g2_fill_1 FILLER_21_421 ();
 sg13g2_decap_4 FILLER_21_427 ();
 sg13g2_fill_2 FILLER_21_431 ();
 sg13g2_fill_2 FILLER_21_455 ();
 sg13g2_fill_2 FILLER_21_460 ();
 sg13g2_decap_4 FILLER_21_467 ();
 sg13g2_fill_1 FILLER_21_471 ();
 sg13g2_fill_2 FILLER_21_486 ();
 sg13g2_fill_2 FILLER_21_496 ();
 sg13g2_fill_2 FILLER_21_526 ();
 sg13g2_decap_8 FILLER_21_547 ();
 sg13g2_fill_2 FILLER_21_567 ();
 sg13g2_fill_1 FILLER_21_569 ();
 sg13g2_decap_4 FILLER_21_575 ();
 sg13g2_fill_1 FILLER_21_579 ();
 sg13g2_decap_8 FILLER_21_626 ();
 sg13g2_decap_4 FILLER_21_633 ();
 sg13g2_fill_2 FILLER_21_637 ();
 sg13g2_fill_2 FILLER_21_648 ();
 sg13g2_fill_1 FILLER_21_650 ();
 sg13g2_decap_8 FILLER_21_682 ();
 sg13g2_decap_8 FILLER_21_689 ();
 sg13g2_fill_2 FILLER_21_696 ();
 sg13g2_decap_4 FILLER_21_703 ();
 sg13g2_fill_2 FILLER_21_707 ();
 sg13g2_decap_4 FILLER_21_760 ();
 sg13g2_fill_1 FILLER_21_764 ();
 sg13g2_fill_2 FILLER_21_821 ();
 sg13g2_fill_1 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_846 ();
 sg13g2_decap_4 FILLER_21_853 ();
 sg13g2_fill_2 FILLER_21_857 ();
 sg13g2_fill_2 FILLER_21_868 ();
 sg13g2_decap_8 FILLER_21_888 ();
 sg13g2_fill_2 FILLER_21_895 ();
 sg13g2_fill_1 FILLER_21_897 ();
 sg13g2_fill_1 FILLER_21_919 ();
 sg13g2_decap_8 FILLER_21_925 ();
 sg13g2_fill_2 FILLER_21_932 ();
 sg13g2_fill_1 FILLER_21_954 ();
 sg13g2_decap_8 FILLER_21_1012 ();
 sg13g2_decap_4 FILLER_21_1019 ();
 sg13g2_fill_2 FILLER_21_1023 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_87 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_decap_4 FILLER_22_113 ();
 sg13g2_decap_8 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_145 ();
 sg13g2_decap_4 FILLER_22_151 ();
 sg13g2_fill_1 FILLER_22_155 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_decap_4 FILLER_22_169 ();
 sg13g2_fill_2 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_261 ();
 sg13g2_decap_8 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_282 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_4 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_416 ();
 sg13g2_fill_1 FILLER_22_423 ();
 sg13g2_decap_8 FILLER_22_430 ();
 sg13g2_decap_8 FILLER_22_437 ();
 sg13g2_fill_2 FILLER_22_444 ();
 sg13g2_fill_1 FILLER_22_446 ();
 sg13g2_fill_1 FILLER_22_461 ();
 sg13g2_fill_2 FILLER_22_477 ();
 sg13g2_fill_2 FILLER_22_539 ();
 sg13g2_fill_1 FILLER_22_592 ();
 sg13g2_fill_2 FILLER_22_654 ();
 sg13g2_decap_8 FILLER_22_692 ();
 sg13g2_decap_8 FILLER_22_699 ();
 sg13g2_fill_1 FILLER_22_727 ();
 sg13g2_fill_1 FILLER_22_745 ();
 sg13g2_decap_8 FILLER_22_755 ();
 sg13g2_decap_4 FILLER_22_762 ();
 sg13g2_fill_2 FILLER_22_766 ();
 sg13g2_fill_2 FILLER_22_794 ();
 sg13g2_decap_8 FILLER_22_832 ();
 sg13g2_decap_8 FILLER_22_839 ();
 sg13g2_decap_4 FILLER_22_890 ();
 sg13g2_decap_8 FILLER_22_902 ();
 sg13g2_fill_1 FILLER_22_909 ();
 sg13g2_decap_8 FILLER_22_914 ();
 sg13g2_fill_1 FILLER_22_921 ();
 sg13g2_fill_2 FILLER_22_944 ();
 sg13g2_decap_8 FILLER_22_955 ();
 sg13g2_decap_4 FILLER_22_962 ();
 sg13g2_fill_2 FILLER_22_979 ();
 sg13g2_decap_4 FILLER_22_985 ();
 sg13g2_fill_2 FILLER_22_989 ();
 sg13g2_decap_8 FILLER_22_1018 ();
 sg13g2_decap_4 FILLER_22_1025 ();
 sg13g2_decap_4 FILLER_23_8 ();
 sg13g2_fill_1 FILLER_23_12 ();
 sg13g2_decap_8 FILLER_23_41 ();
 sg13g2_decap_4 FILLER_23_48 ();
 sg13g2_decap_4 FILLER_23_62 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_decap_4 FILLER_23_131 ();
 sg13g2_fill_2 FILLER_23_146 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_172 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_203 ();
 sg13g2_decap_4 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_253 ();
 sg13g2_decap_8 FILLER_23_260 ();
 sg13g2_decap_8 FILLER_23_267 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_decap_4 FILLER_23_288 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_4 FILLER_23_387 ();
 sg13g2_fill_2 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_4 FILLER_23_455 ();
 sg13g2_fill_1 FILLER_23_459 ();
 sg13g2_decap_8 FILLER_23_471 ();
 sg13g2_decap_4 FILLER_23_482 ();
 sg13g2_fill_2 FILLER_23_491 ();
 sg13g2_fill_1 FILLER_23_493 ();
 sg13g2_fill_2 FILLER_23_510 ();
 sg13g2_fill_2 FILLER_23_533 ();
 sg13g2_fill_1 FILLER_23_535 ();
 sg13g2_fill_2 FILLER_23_541 ();
 sg13g2_decap_4 FILLER_23_637 ();
 sg13g2_fill_1 FILLER_23_641 ();
 sg13g2_fill_2 FILLER_23_650 ();
 sg13g2_decap_8 FILLER_23_670 ();
 sg13g2_fill_2 FILLER_23_677 ();
 sg13g2_fill_2 FILLER_23_729 ();
 sg13g2_fill_1 FILLER_23_731 ();
 sg13g2_fill_2 FILLER_23_741 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_4 FILLER_23_776 ();
 sg13g2_fill_1 FILLER_23_780 ();
 sg13g2_fill_2 FILLER_23_785 ();
 sg13g2_fill_2 FILLER_23_805 ();
 sg13g2_fill_2 FILLER_23_883 ();
 sg13g2_fill_1 FILLER_23_885 ();
 sg13g2_fill_2 FILLER_23_890 ();
 sg13g2_fill_1 FILLER_23_902 ();
 sg13g2_decap_8 FILLER_23_912 ();
 sg13g2_decap_4 FILLER_23_919 ();
 sg13g2_fill_1 FILLER_23_923 ();
 sg13g2_fill_2 FILLER_23_929 ();
 sg13g2_fill_1 FILLER_23_931 ();
 sg13g2_fill_2 FILLER_23_947 ();
 sg13g2_fill_1 FILLER_23_949 ();
 sg13g2_decap_4 FILLER_23_1004 ();
 sg13g2_fill_2 FILLER_23_1008 ();
 sg13g2_decap_8 FILLER_23_1019 ();
 sg13g2_fill_2 FILLER_23_1026 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_4 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_78 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_fill_2 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_decap_4 FILLER_24_237 ();
 sg13g2_fill_2 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_265 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_decap_4 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_4 FILLER_24_327 ();
 sg13g2_decap_4 FILLER_24_342 ();
 sg13g2_fill_2 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_374 ();
 sg13g2_decap_4 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_384 ();
 sg13g2_decap_4 FILLER_24_392 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_401 ();
 sg13g2_fill_2 FILLER_24_405 ();
 sg13g2_fill_2 FILLER_24_425 ();
 sg13g2_fill_2 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_fill_1 FILLER_24_459 ();
 sg13g2_fill_2 FILLER_24_478 ();
 sg13g2_fill_1 FILLER_24_480 ();
 sg13g2_fill_2 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_502 ();
 sg13g2_fill_1 FILLER_24_509 ();
 sg13g2_fill_2 FILLER_24_515 ();
 sg13g2_fill_1 FILLER_24_517 ();
 sg13g2_decap_8 FILLER_24_531 ();
 sg13g2_decap_8 FILLER_24_538 ();
 sg13g2_decap_8 FILLER_24_545 ();
 sg13g2_decap_8 FILLER_24_561 ();
 sg13g2_fill_2 FILLER_24_568 ();
 sg13g2_fill_1 FILLER_24_570 ();
 sg13g2_fill_1 FILLER_24_589 ();
 sg13g2_decap_8 FILLER_24_627 ();
 sg13g2_decap_8 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_641 ();
 sg13g2_fill_2 FILLER_24_648 ();
 sg13g2_decap_8 FILLER_24_670 ();
 sg13g2_decap_8 FILLER_24_677 ();
 sg13g2_fill_2 FILLER_24_688 ();
 sg13g2_fill_1 FILLER_24_690 ();
 sg13g2_fill_2 FILLER_24_766 ();
 sg13g2_fill_1 FILLER_24_777 ();
 sg13g2_fill_1 FILLER_24_783 ();
 sg13g2_fill_2 FILLER_24_820 ();
 sg13g2_fill_1 FILLER_24_822 ();
 sg13g2_fill_1 FILLER_24_877 ();
 sg13g2_fill_2 FILLER_24_890 ();
 sg13g2_fill_1 FILLER_24_892 ();
 sg13g2_decap_4 FILLER_24_924 ();
 sg13g2_fill_1 FILLER_24_928 ();
 sg13g2_fill_1 FILLER_24_942 ();
 sg13g2_fill_2 FILLER_24_954 ();
 sg13g2_decap_8 FILLER_24_968 ();
 sg13g2_decap_8 FILLER_24_975 ();
 sg13g2_decap_8 FILLER_24_982 ();
 sg13g2_decap_8 FILLER_24_989 ();
 sg13g2_decap_8 FILLER_24_996 ();
 sg13g2_decap_8 FILLER_24_1003 ();
 sg13g2_decap_8 FILLER_24_1010 ();
 sg13g2_decap_8 FILLER_24_1017 ();
 sg13g2_decap_4 FILLER_24_1024 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_8 ();
 sg13g2_decap_4 FILLER_25_15 ();
 sg13g2_fill_1 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_75 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_fill_2 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_111 ();
 sg13g2_decap_8 FILLER_25_118 ();
 sg13g2_decap_8 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_180 ();
 sg13g2_fill_1 FILLER_25_182 ();
 sg13g2_decap_4 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_decap_4 FILLER_25_212 ();
 sg13g2_decap_4 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_decap_4 FILLER_25_336 ();
 sg13g2_decap_4 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_348 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_fill_2 FILLER_25_393 ();
 sg13g2_fill_1 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_4 FILLER_25_409 ();
 sg13g2_decap_8 FILLER_25_449 ();
 sg13g2_decap_8 FILLER_25_456 ();
 sg13g2_decap_8 FILLER_25_463 ();
 sg13g2_fill_1 FILLER_25_482 ();
 sg13g2_decap_4 FILLER_25_501 ();
 sg13g2_fill_2 FILLER_25_505 ();
 sg13g2_fill_2 FILLER_25_520 ();
 sg13g2_fill_1 FILLER_25_522 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_fill_1 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_decap_8 FILLER_25_564 ();
 sg13g2_decap_4 FILLER_25_571 ();
 sg13g2_fill_2 FILLER_25_588 ();
 sg13g2_fill_2 FILLER_25_606 ();
 sg13g2_fill_1 FILLER_25_608 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_decap_4 FILLER_25_629 ();
 sg13g2_decap_4 FILLER_25_661 ();
 sg13g2_fill_2 FILLER_25_665 ();
 sg13g2_decap_4 FILLER_25_675 ();
 sg13g2_fill_2 FILLER_25_679 ();
 sg13g2_decap_4 FILLER_25_685 ();
 sg13g2_fill_1 FILLER_25_689 ();
 sg13g2_fill_1 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_734 ();
 sg13g2_fill_2 FILLER_25_741 ();
 sg13g2_fill_1 FILLER_25_787 ();
 sg13g2_decap_8 FILLER_25_820 ();
 sg13g2_decap_8 FILLER_25_827 ();
 sg13g2_decap_4 FILLER_25_834 ();
 sg13g2_fill_2 FILLER_25_838 ();
 sg13g2_decap_8 FILLER_25_862 ();
 sg13g2_decap_8 FILLER_25_869 ();
 sg13g2_decap_8 FILLER_25_876 ();
 sg13g2_decap_4 FILLER_25_883 ();
 sg13g2_fill_1 FILLER_25_887 ();
 sg13g2_fill_1 FILLER_25_933 ();
 sg13g2_fill_2 FILLER_25_938 ();
 sg13g2_decap_8 FILLER_25_958 ();
 sg13g2_decap_4 FILLER_25_965 ();
 sg13g2_fill_1 FILLER_25_969 ();
 sg13g2_decap_8 FILLER_25_998 ();
 sg13g2_decap_8 FILLER_25_1005 ();
 sg13g2_decap_8 FILLER_25_1012 ();
 sg13g2_decap_8 FILLER_25_1019 ();
 sg13g2_fill_2 FILLER_25_1026 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_39 ();
 sg13g2_fill_2 FILLER_26_43 ();
 sg13g2_fill_1 FILLER_26_90 ();
 sg13g2_decap_4 FILLER_26_101 ();
 sg13g2_fill_2 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_127 ();
 sg13g2_decap_4 FILLER_26_134 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_4 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_171 ();
 sg13g2_decap_4 FILLER_26_188 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_8 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_4 FILLER_26_375 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_412 ();
 sg13g2_fill_2 FILLER_26_419 ();
 sg13g2_fill_1 FILLER_26_421 ();
 sg13g2_decap_8 FILLER_26_425 ();
 sg13g2_fill_2 FILLER_26_432 ();
 sg13g2_fill_1 FILLER_26_434 ();
 sg13g2_fill_2 FILLER_26_464 ();
 sg13g2_fill_2 FILLER_26_475 ();
 sg13g2_fill_1 FILLER_26_477 ();
 sg13g2_decap_4 FILLER_26_534 ();
 sg13g2_fill_1 FILLER_26_538 ();
 sg13g2_decap_8 FILLER_26_544 ();
 sg13g2_fill_1 FILLER_26_597 ();
 sg13g2_decap_8 FILLER_26_615 ();
 sg13g2_decap_8 FILLER_26_627 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_fill_1 FILLER_26_651 ();
 sg13g2_fill_2 FILLER_26_657 ();
 sg13g2_fill_1 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_699 ();
 sg13g2_decap_8 FILLER_26_706 ();
 sg13g2_decap_8 FILLER_26_713 ();
 sg13g2_decap_8 FILLER_26_720 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_fill_1 FILLER_26_747 ();
 sg13g2_fill_2 FILLER_26_757 ();
 sg13g2_fill_1 FILLER_26_759 ();
 sg13g2_fill_2 FILLER_26_774 ();
 sg13g2_fill_1 FILLER_26_776 ();
 sg13g2_fill_2 FILLER_26_804 ();
 sg13g2_fill_1 FILLER_26_806 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_4 FILLER_26_831 ();
 sg13g2_fill_2 FILLER_26_848 ();
 sg13g2_decap_4 FILLER_26_878 ();
 sg13g2_fill_2 FILLER_26_888 ();
 sg13g2_fill_1 FILLER_26_890 ();
 sg13g2_fill_2 FILLER_26_897 ();
 sg13g2_fill_1 FILLER_26_930 ();
 sg13g2_fill_1 FILLER_26_940 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_decap_8 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_1001 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_decap_4 FILLER_27_16 ();
 sg13g2_decap_8 FILLER_27_38 ();
 sg13g2_decap_8 FILLER_27_58 ();
 sg13g2_fill_1 FILLER_27_93 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_206 ();
 sg13g2_decap_4 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_decap_4 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_decap_4 FILLER_27_293 ();
 sg13g2_fill_2 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_304 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_fill_2 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_366 ();
 sg13g2_decap_4 FILLER_27_373 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_decap_4 FILLER_27_383 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_decap_8 FILLER_27_458 ();
 sg13g2_decap_4 FILLER_27_465 ();
 sg13g2_decap_8 FILLER_27_495 ();
 sg13g2_decap_8 FILLER_27_502 ();
 sg13g2_decap_4 FILLER_27_509 ();
 sg13g2_fill_1 FILLER_27_519 ();
 sg13g2_fill_2 FILLER_27_529 ();
 sg13g2_fill_1 FILLER_27_531 ();
 sg13g2_fill_2 FILLER_27_567 ();
 sg13g2_fill_1 FILLER_27_605 ();
 sg13g2_decap_4 FILLER_27_627 ();
 sg13g2_fill_1 FILLER_27_631 ();
 sg13g2_decap_4 FILLER_27_638 ();
 sg13g2_fill_1 FILLER_27_642 ();
 sg13g2_fill_1 FILLER_27_654 ();
 sg13g2_decap_4 FILLER_27_686 ();
 sg13g2_fill_2 FILLER_27_729 ();
 sg13g2_fill_2 FILLER_27_803 ();
 sg13g2_fill_2 FILLER_27_827 ();
 sg13g2_fill_1 FILLER_27_860 ();
 sg13g2_decap_4 FILLER_27_876 ();
 sg13g2_decap_4 FILLER_27_884 ();
 sg13g2_fill_2 FILLER_27_888 ();
 sg13g2_decap_4 FILLER_27_898 ();
 sg13g2_fill_2 FILLER_27_902 ();
 sg13g2_fill_1 FILLER_27_909 ();
 sg13g2_decap_8 FILLER_27_976 ();
 sg13g2_fill_2 FILLER_27_983 ();
 sg13g2_fill_1 FILLER_27_985 ();
 sg13g2_decap_8 FILLER_27_999 ();
 sg13g2_decap_8 FILLER_27_1006 ();
 sg13g2_decap_8 FILLER_27_1013 ();
 sg13g2_decap_8 FILLER_27_1020 ();
 sg13g2_fill_2 FILLER_27_1027 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_33 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_4 FILLER_28_84 ();
 sg13g2_fill_1 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_decap_4 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_decap_4 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_301 ();
 sg13g2_decap_4 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_331 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_fill_2 FILLER_28_358 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_387 ();
 sg13g2_fill_1 FILLER_28_397 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_fill_2 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_440 ();
 sg13g2_decap_4 FILLER_28_448 ();
 sg13g2_decap_4 FILLER_28_489 ();
 sg13g2_fill_2 FILLER_28_493 ();
 sg13g2_decap_4 FILLER_28_499 ();
 sg13g2_fill_2 FILLER_28_503 ();
 sg13g2_decap_8 FILLER_28_524 ();
 sg13g2_fill_2 FILLER_28_531 ();
 sg13g2_fill_1 FILLER_28_533 ();
 sg13g2_decap_8 FILLER_28_543 ();
 sg13g2_decap_4 FILLER_28_550 ();
 sg13g2_fill_1 FILLER_28_567 ();
 sg13g2_decap_4 FILLER_28_596 ();
 sg13g2_fill_1 FILLER_28_620 ();
 sg13g2_decap_4 FILLER_28_624 ();
 sg13g2_decap_4 FILLER_28_634 ();
 sg13g2_fill_1 FILLER_28_638 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_fill_2 FILLER_28_666 ();
 sg13g2_fill_2 FILLER_28_691 ();
 sg13g2_fill_2 FILLER_28_707 ();
 sg13g2_fill_2 FILLER_28_716 ();
 sg13g2_fill_2 FILLER_28_736 ();
 sg13g2_fill_2 FILLER_28_774 ();
 sg13g2_fill_1 FILLER_28_776 ();
 sg13g2_decap_4 FILLER_28_799 ();
 sg13g2_fill_1 FILLER_28_803 ();
 sg13g2_decap_4 FILLER_28_832 ();
 sg13g2_fill_1 FILLER_28_836 ();
 sg13g2_fill_2 FILLER_28_846 ();
 sg13g2_fill_1 FILLER_28_860 ();
 sg13g2_fill_2 FILLER_28_891 ();
 sg13g2_decap_8 FILLER_28_897 ();
 sg13g2_decap_4 FILLER_28_904 ();
 sg13g2_fill_1 FILLER_28_908 ();
 sg13g2_decap_8 FILLER_28_914 ();
 sg13g2_fill_2 FILLER_28_921 ();
 sg13g2_fill_1 FILLER_28_929 ();
 sg13g2_decap_8 FILLER_28_956 ();
 sg13g2_decap_8 FILLER_28_963 ();
 sg13g2_decap_8 FILLER_28_970 ();
 sg13g2_decap_8 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_984 ();
 sg13g2_decap_8 FILLER_28_991 ();
 sg13g2_decap_8 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1005 ();
 sg13g2_decap_8 FILLER_28_1012 ();
 sg13g2_decap_8 FILLER_28_1019 ();
 sg13g2_fill_2 FILLER_28_1026 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_fill_2 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_16 ();
 sg13g2_fill_2 FILLER_29_23 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_fill_2 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_61 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_decap_4 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_fill_1 FILLER_29_179 ();
 sg13g2_fill_1 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_decap_4 FILLER_29_230 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_265 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_294 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_4 FILLER_29_364 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_decap_4 FILLER_29_401 ();
 sg13g2_decap_4 FILLER_29_410 ();
 sg13g2_fill_1 FILLER_29_414 ();
 sg13g2_decap_4 FILLER_29_420 ();
 sg13g2_fill_1 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_478 ();
 sg13g2_decap_4 FILLER_29_507 ();
 sg13g2_fill_1 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_fill_2 FILLER_29_545 ();
 sg13g2_fill_1 FILLER_29_547 ();
 sg13g2_fill_2 FILLER_29_567 ();
 sg13g2_fill_2 FILLER_29_616 ();
 sg13g2_fill_1 FILLER_29_618 ();
 sg13g2_decap_8 FILLER_29_624 ();
 sg13g2_decap_8 FILLER_29_631 ();
 sg13g2_fill_2 FILLER_29_638 ();
 sg13g2_fill_1 FILLER_29_640 ();
 sg13g2_fill_2 FILLER_29_656 ();
 sg13g2_fill_2 FILLER_29_665 ();
 sg13g2_fill_1 FILLER_29_671 ();
 sg13g2_decap_4 FILLER_29_687 ();
 sg13g2_fill_1 FILLER_29_691 ();
 sg13g2_decap_4 FILLER_29_696 ();
 sg13g2_fill_1 FILLER_29_700 ();
 sg13g2_fill_2 FILLER_29_709 ();
 sg13g2_fill_1 FILLER_29_726 ();
 sg13g2_fill_1 FILLER_29_736 ();
 sg13g2_decap_8 FILLER_29_764 ();
 sg13g2_fill_2 FILLER_29_771 ();
 sg13g2_fill_2 FILLER_29_777 ();
 sg13g2_fill_1 FILLER_29_779 ();
 sg13g2_fill_2 FILLER_29_799 ();
 sg13g2_decap_4 FILLER_29_815 ();
 sg13g2_fill_1 FILLER_29_819 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_decap_8 FILLER_29_901 ();
 sg13g2_decap_4 FILLER_29_908 ();
 sg13g2_fill_2 FILLER_29_912 ();
 sg13g2_decap_8 FILLER_29_958 ();
 sg13g2_decap_8 FILLER_29_965 ();
 sg13g2_decap_8 FILLER_29_972 ();
 sg13g2_decap_8 FILLER_29_979 ();
 sg13g2_decap_8 FILLER_29_986 ();
 sg13g2_decap_8 FILLER_29_993 ();
 sg13g2_decap_8 FILLER_29_1000 ();
 sg13g2_decap_8 FILLER_29_1007 ();
 sg13g2_decap_8 FILLER_29_1014 ();
 sg13g2_decap_8 FILLER_29_1021 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_6 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_decap_8 FILLER_30_54 ();
 sg13g2_decap_4 FILLER_30_61 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_fill_2 FILLER_30_94 ();
 sg13g2_decap_4 FILLER_30_124 ();
 sg13g2_decap_8 FILLER_30_174 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_fill_2 FILLER_30_272 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_331 ();
 sg13g2_fill_1 FILLER_30_333 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_365 ();
 sg13g2_decap_4 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_385 ();
 sg13g2_fill_1 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_8 FILLER_30_424 ();
 sg13g2_decap_8 FILLER_30_431 ();
 sg13g2_fill_1 FILLER_30_468 ();
 sg13g2_fill_2 FILLER_30_487 ();
 sg13g2_fill_2 FILLER_30_526 ();
 sg13g2_fill_1 FILLER_30_528 ();
 sg13g2_decap_8 FILLER_30_557 ();
 sg13g2_decap_8 FILLER_30_564 ();
 sg13g2_decap_4 FILLER_30_571 ();
 sg13g2_fill_2 FILLER_30_575 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_4 FILLER_30_588 ();
 sg13g2_fill_1 FILLER_30_592 ();
 sg13g2_fill_1 FILLER_30_612 ();
 sg13g2_fill_2 FILLER_30_629 ();
 sg13g2_decap_4 FILLER_30_635 ();
 sg13g2_fill_2 FILLER_30_639 ();
 sg13g2_fill_2 FILLER_30_652 ();
 sg13g2_fill_1 FILLER_30_654 ();
 sg13g2_fill_2 FILLER_30_660 ();
 sg13g2_fill_1 FILLER_30_662 ();
 sg13g2_decap_4 FILLER_30_685 ();
 sg13g2_fill_2 FILLER_30_689 ();
 sg13g2_fill_2 FILLER_30_700 ();
 sg13g2_fill_2 FILLER_30_726 ();
 sg13g2_fill_1 FILLER_30_735 ();
 sg13g2_decap_4 FILLER_30_763 ();
 sg13g2_fill_1 FILLER_30_767 ();
 sg13g2_decap_4 FILLER_30_796 ();
 sg13g2_fill_2 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_fill_2 FILLER_30_852 ();
 sg13g2_fill_1 FILLER_30_854 ();
 sg13g2_fill_2 FILLER_30_920 ();
 sg13g2_decap_8 FILLER_30_949 ();
 sg13g2_decap_8 FILLER_30_956 ();
 sg13g2_decap_8 FILLER_30_963 ();
 sg13g2_decap_8 FILLER_30_970 ();
 sg13g2_decap_8 FILLER_30_977 ();
 sg13g2_decap_8 FILLER_30_984 ();
 sg13g2_decap_8 FILLER_30_991 ();
 sg13g2_decap_8 FILLER_30_998 ();
 sg13g2_decap_8 FILLER_30_1005 ();
 sg13g2_decap_8 FILLER_30_1012 ();
 sg13g2_decap_4 FILLER_30_1019 ();
 sg13g2_fill_2 FILLER_30_1023 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_decap_4 FILLER_31_16 ();
 sg13g2_fill_2 FILLER_31_20 ();
 sg13g2_decap_4 FILLER_31_31 ();
 sg13g2_decap_4 FILLER_31_83 ();
 sg13g2_fill_2 FILLER_31_87 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_fill_2 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_decap_8 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_242 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_4 FILLER_31_273 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_decap_4 FILLER_31_369 ();
 sg13g2_fill_2 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_fill_2 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_403 ();
 sg13g2_decap_8 FILLER_31_410 ();
 sg13g2_decap_8 FILLER_31_417 ();
 sg13g2_fill_2 FILLER_31_424 ();
 sg13g2_decap_8 FILLER_31_431 ();
 sg13g2_decap_8 FILLER_31_438 ();
 sg13g2_fill_2 FILLER_31_445 ();
 sg13g2_fill_1 FILLER_31_447 ();
 sg13g2_fill_2 FILLER_31_485 ();
 sg13g2_decap_8 FILLER_31_500 ();
 sg13g2_decap_8 FILLER_31_507 ();
 sg13g2_decap_8 FILLER_31_514 ();
 sg13g2_decap_8 FILLER_31_521 ();
 sg13g2_decap_4 FILLER_31_528 ();
 sg13g2_fill_1 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_538 ();
 sg13g2_decap_8 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_552 ();
 sg13g2_decap_8 FILLER_31_587 ();
 sg13g2_decap_8 FILLER_31_613 ();
 sg13g2_decap_4 FILLER_31_646 ();
 sg13g2_fill_1 FILLER_31_650 ();
 sg13g2_decap_4 FILLER_31_655 ();
 sg13g2_fill_1 FILLER_31_659 ();
 sg13g2_fill_1 FILLER_31_664 ();
 sg13g2_fill_2 FILLER_31_701 ();
 sg13g2_fill_1 FILLER_31_703 ();
 sg13g2_fill_1 FILLER_31_713 ();
 sg13g2_fill_2 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_4 FILLER_31_784 ();
 sg13g2_fill_1 FILLER_31_788 ();
 sg13g2_decap_4 FILLER_31_816 ();
 sg13g2_fill_1 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_831 ();
 sg13g2_fill_2 FILLER_31_838 ();
 sg13g2_decap_4 FILLER_31_846 ();
 sg13g2_fill_2 FILLER_31_850 ();
 sg13g2_fill_2 FILLER_31_874 ();
 sg13g2_fill_1 FILLER_31_876 ();
 sg13g2_fill_1 FILLER_31_887 ();
 sg13g2_fill_1 FILLER_31_906 ();
 sg13g2_fill_1 FILLER_31_916 ();
 sg13g2_decap_8 FILLER_31_954 ();
 sg13g2_decap_8 FILLER_31_961 ();
 sg13g2_decap_8 FILLER_31_968 ();
 sg13g2_decap_8 FILLER_31_975 ();
 sg13g2_decap_8 FILLER_31_982 ();
 sg13g2_decap_8 FILLER_31_989 ();
 sg13g2_decap_8 FILLER_31_996 ();
 sg13g2_decap_8 FILLER_31_1003 ();
 sg13g2_decap_8 FILLER_31_1010 ();
 sg13g2_decap_8 FILLER_31_1017 ();
 sg13g2_decap_4 FILLER_31_1024 ();
 sg13g2_fill_1 FILLER_31_1028 ();
 sg13g2_decap_4 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_8 ();
 sg13g2_decap_4 FILLER_32_37 ();
 sg13g2_fill_2 FILLER_32_41 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_decap_4 FILLER_32_178 ();
 sg13g2_decap_4 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_385 ();
 sg13g2_fill_2 FILLER_32_395 ();
 sg13g2_fill_2 FILLER_32_403 ();
 sg13g2_fill_1 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_32_411 ();
 sg13g2_fill_1 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_4 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_456 ();
 sg13g2_fill_2 FILLER_32_463 ();
 sg13g2_fill_1 FILLER_32_487 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_4 FILLER_32_518 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_decap_8 FILLER_32_548 ();
 sg13g2_fill_2 FILLER_32_555 ();
 sg13g2_fill_1 FILLER_32_557 ();
 sg13g2_fill_2 FILLER_32_577 ();
 sg13g2_fill_1 FILLER_32_579 ();
 sg13g2_decap_8 FILLER_32_589 ();
 sg13g2_decap_4 FILLER_32_596 ();
 sg13g2_decap_4 FILLER_32_624 ();
 sg13g2_fill_2 FILLER_32_628 ();
 sg13g2_decap_8 FILLER_32_652 ();
 sg13g2_fill_2 FILLER_32_659 ();
 sg13g2_fill_1 FILLER_32_679 ();
 sg13g2_decap_4 FILLER_32_693 ();
 sg13g2_fill_2 FILLER_32_697 ();
 sg13g2_fill_2 FILLER_32_776 ();
 sg13g2_decap_4 FILLER_32_852 ();
 sg13g2_fill_2 FILLER_32_856 ();
 sg13g2_fill_1 FILLER_32_896 ();
 sg13g2_decap_8 FILLER_32_943 ();
 sg13g2_decap_8 FILLER_32_950 ();
 sg13g2_decap_8 FILLER_32_957 ();
 sg13g2_decap_8 FILLER_32_964 ();
 sg13g2_decap_8 FILLER_32_971 ();
 sg13g2_decap_8 FILLER_32_978 ();
 sg13g2_decap_8 FILLER_32_985 ();
 sg13g2_decap_8 FILLER_32_992 ();
 sg13g2_decap_8 FILLER_32_999 ();
 sg13g2_decap_8 FILLER_32_1006 ();
 sg13g2_decap_8 FILLER_32_1013 ();
 sg13g2_decap_8 FILLER_32_1020 ();
 sg13g2_fill_2 FILLER_32_1027 ();
 sg13g2_decap_8 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_decap_4 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_22 ();
 sg13g2_decap_8 FILLER_33_32 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_4 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_decap_4 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_4 FILLER_33_387 ();
 sg13g2_decap_4 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_33_440 ();
 sg13g2_fill_1 FILLER_33_478 ();
 sg13g2_decap_8 FILLER_33_516 ();
 sg13g2_decap_4 FILLER_33_528 ();
 sg13g2_decap_8 FILLER_33_545 ();
 sg13g2_decap_4 FILLER_33_552 ();
 sg13g2_decap_4 FILLER_33_597 ();
 sg13g2_fill_1 FILLER_33_601 ();
 sg13g2_decap_4 FILLER_33_618 ();
 sg13g2_fill_1 FILLER_33_622 ();
 sg13g2_fill_2 FILLER_33_633 ();
 sg13g2_fill_1 FILLER_33_644 ();
 sg13g2_fill_1 FILLER_33_673 ();
 sg13g2_fill_1 FILLER_33_687 ();
 sg13g2_decap_8 FILLER_33_758 ();
 sg13g2_decap_4 FILLER_33_765 ();
 sg13g2_decap_4 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_837 ();
 sg13g2_decap_8 FILLER_33_844 ();
 sg13g2_fill_2 FILLER_33_851 ();
 sg13g2_fill_1 FILLER_33_853 ();
 sg13g2_decap_8 FILLER_33_873 ();
 sg13g2_fill_2 FILLER_33_880 ();
 sg13g2_fill_1 FILLER_33_882 ();
 sg13g2_decap_4 FILLER_33_911 ();
 sg13g2_fill_1 FILLER_33_915 ();
 sg13g2_decap_8 FILLER_33_944 ();
 sg13g2_decap_8 FILLER_33_951 ();
 sg13g2_decap_8 FILLER_33_958 ();
 sg13g2_decap_8 FILLER_33_965 ();
 sg13g2_decap_8 FILLER_33_972 ();
 sg13g2_decap_8 FILLER_33_979 ();
 sg13g2_decap_8 FILLER_33_986 ();
 sg13g2_decap_8 FILLER_33_993 ();
 sg13g2_decap_8 FILLER_33_1000 ();
 sg13g2_decap_8 FILLER_33_1007 ();
 sg13g2_decap_8 FILLER_33_1014 ();
 sg13g2_decap_8 FILLER_33_1021 ();
 sg13g2_fill_1 FILLER_33_1028 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_2 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_decap_4 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_decap_4 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_decap_4 FILLER_34_394 ();
 sg13g2_fill_1 FILLER_34_398 ();
 sg13g2_decap_8 FILLER_34_407 ();
 sg13g2_decap_4 FILLER_34_414 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_decap_8 FILLER_34_430 ();
 sg13g2_decap_8 FILLER_34_437 ();
 sg13g2_decap_4 FILLER_34_444 ();
 sg13g2_fill_1 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_456 ();
 sg13g2_fill_1 FILLER_34_463 ();
 sg13g2_fill_1 FILLER_34_492 ();
 sg13g2_decap_4 FILLER_34_499 ();
 sg13g2_fill_1 FILLER_34_530 ();
 sg13g2_fill_2 FILLER_34_559 ();
 sg13g2_fill_2 FILLER_34_584 ();
 sg13g2_fill_1 FILLER_34_586 ();
 sg13g2_decap_8 FILLER_34_596 ();
 sg13g2_fill_1 FILLER_34_603 ();
 sg13g2_fill_1 FILLER_34_697 ();
 sg13g2_decap_4 FILLER_34_712 ();
 sg13g2_fill_2 FILLER_34_729 ();
 sg13g2_decap_4 FILLER_34_736 ();
 sg13g2_fill_1 FILLER_34_740 ();
 sg13g2_decap_8 FILLER_34_759 ();
 sg13g2_decap_8 FILLER_34_766 ();
 sg13g2_fill_2 FILLER_34_773 ();
 sg13g2_fill_1 FILLER_34_775 ();
 sg13g2_fill_2 FILLER_34_789 ();
 sg13g2_decap_4 FILLER_34_836 ();
 sg13g2_fill_1 FILLER_34_840 ();
 sg13g2_decap_4 FILLER_34_868 ();
 sg13g2_fill_1 FILLER_34_872 ();
 sg13g2_fill_2 FILLER_34_877 ();
 sg13g2_fill_2 FILLER_34_892 ();
 sg13g2_fill_1 FILLER_34_894 ();
 sg13g2_decap_4 FILLER_34_899 ();
 sg13g2_fill_1 FILLER_34_920 ();
 sg13g2_decap_8 FILLER_34_924 ();
 sg13g2_decap_8 FILLER_34_931 ();
 sg13g2_decap_8 FILLER_34_938 ();
 sg13g2_decap_8 FILLER_34_945 ();
 sg13g2_decap_8 FILLER_34_952 ();
 sg13g2_decap_8 FILLER_34_959 ();
 sg13g2_decap_8 FILLER_34_966 ();
 sg13g2_decap_8 FILLER_34_973 ();
 sg13g2_decap_8 FILLER_34_980 ();
 sg13g2_decap_8 FILLER_34_987 ();
 sg13g2_decap_8 FILLER_34_994 ();
 sg13g2_decap_8 FILLER_34_1001 ();
 sg13g2_decap_8 FILLER_34_1008 ();
 sg13g2_decap_8 FILLER_34_1015 ();
 sg13g2_decap_8 FILLER_34_1022 ();
 sg13g2_decap_8 FILLER_35_41 ();
 sg13g2_fill_2 FILLER_35_48 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_decap_4 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_203 ();
 sg13g2_decap_4 FILLER_35_223 ();
 sg13g2_decap_4 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_decap_8 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_272 ();
 sg13g2_decap_4 FILLER_35_283 ();
 sg13g2_decap_4 FILLER_35_324 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_decap_4 FILLER_35_380 ();
 sg13g2_decap_4 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_426 ();
 sg13g2_fill_2 FILLER_35_433 ();
 sg13g2_fill_1 FILLER_35_448 ();
 sg13g2_fill_2 FILLER_35_486 ();
 sg13g2_fill_2 FILLER_35_518 ();
 sg13g2_fill_1 FILLER_35_520 ();
 sg13g2_fill_2 FILLER_35_538 ();
 sg13g2_fill_1 FILLER_35_540 ();
 sg13g2_decap_4 FILLER_35_545 ();
 sg13g2_fill_2 FILLER_35_549 ();
 sg13g2_decap_8 FILLER_35_597 ();
 sg13g2_fill_2 FILLER_35_604 ();
 sg13g2_fill_1 FILLER_35_606 ();
 sg13g2_fill_2 FILLER_35_617 ();
 sg13g2_decap_8 FILLER_35_624 ();
 sg13g2_decap_4 FILLER_35_631 ();
 sg13g2_fill_1 FILLER_35_639 ();
 sg13g2_fill_1 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_fill_2 FILLER_35_693 ();
 sg13g2_fill_1 FILLER_35_695 ();
 sg13g2_decap_4 FILLER_35_728 ();
 sg13g2_decap_4 FILLER_35_758 ();
 sg13g2_fill_1 FILLER_35_790 ();
 sg13g2_fill_2 FILLER_35_819 ();
 sg13g2_fill_1 FILLER_35_821 ();
 sg13g2_fill_1 FILLER_35_835 ();
 sg13g2_fill_1 FILLER_35_859 ();
 sg13g2_fill_2 FILLER_35_873 ();
 sg13g2_decap_8 FILLER_35_936 ();
 sg13g2_decap_8 FILLER_35_943 ();
 sg13g2_decap_8 FILLER_35_950 ();
 sg13g2_decap_8 FILLER_35_957 ();
 sg13g2_decap_8 FILLER_35_964 ();
 sg13g2_decap_8 FILLER_35_971 ();
 sg13g2_decap_8 FILLER_35_978 ();
 sg13g2_decap_8 FILLER_35_985 ();
 sg13g2_decap_8 FILLER_35_992 ();
 sg13g2_decap_8 FILLER_35_999 ();
 sg13g2_decap_8 FILLER_35_1006 ();
 sg13g2_decap_8 FILLER_35_1013 ();
 sg13g2_decap_8 FILLER_35_1020 ();
 sg13g2_fill_2 FILLER_35_1027 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_decap_4 FILLER_36_16 ();
 sg13g2_decap_8 FILLER_36_93 ();
 sg13g2_decap_8 FILLER_36_136 ();
 sg13g2_decap_4 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_412 ();
 sg13g2_fill_2 FILLER_36_419 ();
 sg13g2_fill_2 FILLER_36_438 ();
 sg13g2_fill_1 FILLER_36_440 ();
 sg13g2_decap_8 FILLER_36_447 ();
 sg13g2_fill_2 FILLER_36_454 ();
 sg13g2_decap_8 FILLER_36_460 ();
 sg13g2_decap_8 FILLER_36_467 ();
 sg13g2_decap_8 FILLER_36_474 ();
 sg13g2_fill_2 FILLER_36_503 ();
 sg13g2_fill_1 FILLER_36_505 ();
 sg13g2_fill_1 FILLER_36_515 ();
 sg13g2_fill_2 FILLER_36_521 ();
 sg13g2_fill_1 FILLER_36_523 ();
 sg13g2_decap_4 FILLER_36_540 ();
 sg13g2_fill_2 FILLER_36_544 ();
 sg13g2_decap_8 FILLER_36_557 ();
 sg13g2_decap_8 FILLER_36_564 ();
 sg13g2_fill_2 FILLER_36_571 ();
 sg13g2_fill_1 FILLER_36_573 ();
 sg13g2_fill_2 FILLER_36_615 ();
 sg13g2_fill_2 FILLER_36_631 ();
 sg13g2_fill_1 FILLER_36_633 ();
 sg13g2_fill_2 FILLER_36_639 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_fill_2 FILLER_36_665 ();
 sg13g2_fill_1 FILLER_36_667 ();
 sg13g2_decap_8 FILLER_36_696 ();
 sg13g2_decap_4 FILLER_36_703 ();
 sg13g2_decap_8 FILLER_36_724 ();
 sg13g2_decap_4 FILLER_36_731 ();
 sg13g2_fill_1 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_753 ();
 sg13g2_decap_4 FILLER_36_760 ();
 sg13g2_fill_1 FILLER_36_764 ();
 sg13g2_fill_2 FILLER_36_798 ();
 sg13g2_fill_2 FILLER_36_814 ();
 sg13g2_fill_2 FILLER_36_830 ();
 sg13g2_fill_1 FILLER_36_864 ();
 sg13g2_fill_1 FILLER_36_879 ();
 sg13g2_fill_2 FILLER_36_889 ();
 sg13g2_fill_2 FILLER_36_908 ();
 sg13g2_decap_8 FILLER_36_933 ();
 sg13g2_decap_8 FILLER_36_940 ();
 sg13g2_decap_8 FILLER_36_947 ();
 sg13g2_decap_8 FILLER_36_954 ();
 sg13g2_decap_8 FILLER_36_961 ();
 sg13g2_decap_8 FILLER_36_968 ();
 sg13g2_decap_8 FILLER_36_975 ();
 sg13g2_decap_8 FILLER_36_982 ();
 sg13g2_decap_8 FILLER_36_989 ();
 sg13g2_decap_8 FILLER_36_996 ();
 sg13g2_decap_8 FILLER_36_1003 ();
 sg13g2_decap_8 FILLER_36_1010 ();
 sg13g2_decap_8 FILLER_36_1017 ();
 sg13g2_decap_4 FILLER_36_1024 ();
 sg13g2_fill_1 FILLER_36_1028 ();
 sg13g2_decap_4 FILLER_37_27 ();
 sg13g2_fill_2 FILLER_37_31 ();
 sg13g2_fill_1 FILLER_37_75 ();
 sg13g2_decap_8 FILLER_37_89 ();
 sg13g2_decap_8 FILLER_37_96 ();
 sg13g2_decap_4 FILLER_37_103 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_fill_1 FILLER_37_153 ();
 sg13g2_fill_1 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_4 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_207 ();
 sg13g2_fill_2 FILLER_37_222 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_293 ();
 sg13g2_decap_8 FILLER_37_300 ();
 sg13g2_decap_8 FILLER_37_307 ();
 sg13g2_decap_8 FILLER_37_314 ();
 sg13g2_decap_4 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_decap_4 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_2 FILLER_37_418 ();
 sg13g2_decap_8 FILLER_37_443 ();
 sg13g2_fill_1 FILLER_37_450 ();
 sg13g2_fill_2 FILLER_37_456 ();
 sg13g2_decap_8 FILLER_37_464 ();
 sg13g2_decap_8 FILLER_37_471 ();
 sg13g2_fill_2 FILLER_37_478 ();
 sg13g2_fill_1 FILLER_37_480 ();
 sg13g2_fill_2 FILLER_37_490 ();
 sg13g2_fill_2 FILLER_37_510 ();
 sg13g2_fill_1 FILLER_37_527 ();
 sg13g2_decap_4 FILLER_37_536 ();
 sg13g2_fill_2 FILLER_37_540 ();
 sg13g2_fill_2 FILLER_37_550 ();
 sg13g2_fill_1 FILLER_37_552 ();
 sg13g2_decap_8 FILLER_37_571 ();
 sg13g2_decap_8 FILLER_37_578 ();
 sg13g2_decap_4 FILLER_37_585 ();
 sg13g2_fill_2 FILLER_37_589 ();
 sg13g2_fill_1 FILLER_37_600 ();
 sg13g2_fill_1 FILLER_37_624 ();
 sg13g2_decap_4 FILLER_37_638 ();
 sg13g2_fill_1 FILLER_37_642 ();
 sg13g2_decap_8 FILLER_37_656 ();
 sg13g2_decap_8 FILLER_37_663 ();
 sg13g2_decap_8 FILLER_37_670 ();
 sg13g2_decap_4 FILLER_37_677 ();
 sg13g2_fill_2 FILLER_37_681 ();
 sg13g2_decap_4 FILLER_37_711 ();
 sg13g2_fill_1 FILLER_37_715 ();
 sg13g2_decap_8 FILLER_37_724 ();
 sg13g2_decap_8 FILLER_37_731 ();
 sg13g2_decap_8 FILLER_37_761 ();
 sg13g2_decap_8 FILLER_37_768 ();
 sg13g2_fill_2 FILLER_37_775 ();
 sg13g2_fill_1 FILLER_37_777 ();
 sg13g2_fill_1 FILLER_37_791 ();
 sg13g2_fill_1 FILLER_37_815 ();
 sg13g2_fill_2 FILLER_37_832 ();
 sg13g2_fill_1 FILLER_37_853 ();
 sg13g2_decap_4 FILLER_37_882 ();
 sg13g2_fill_1 FILLER_37_886 ();
 sg13g2_decap_8 FILLER_37_926 ();
 sg13g2_decap_8 FILLER_37_933 ();
 sg13g2_decap_8 FILLER_37_940 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_decap_8 FILLER_37_954 ();
 sg13g2_decap_8 FILLER_37_961 ();
 sg13g2_decap_8 FILLER_37_968 ();
 sg13g2_decap_8 FILLER_37_975 ();
 sg13g2_decap_8 FILLER_37_982 ();
 sg13g2_decap_8 FILLER_37_989 ();
 sg13g2_decap_8 FILLER_37_996 ();
 sg13g2_decap_8 FILLER_37_1003 ();
 sg13g2_decap_8 FILLER_37_1010 ();
 sg13g2_decap_8 FILLER_37_1017 ();
 sg13g2_decap_4 FILLER_37_1024 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_decap_8 FILLER_38_128 ();
 sg13g2_decap_4 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_decap_8 FILLER_38_157 ();
 sg13g2_fill_2 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_4 FILLER_38_213 ();
 sg13g2_fill_2 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_fill_2 FILLER_38_411 ();
 sg13g2_fill_1 FILLER_38_413 ();
 sg13g2_fill_2 FILLER_38_424 ();
 sg13g2_fill_1 FILLER_38_426 ();
 sg13g2_decap_4 FILLER_38_441 ();
 sg13g2_fill_2 FILLER_38_445 ();
 sg13g2_decap_8 FILLER_38_464 ();
 sg13g2_decap_8 FILLER_38_471 ();
 sg13g2_fill_1 FILLER_38_478 ();
 sg13g2_fill_2 FILLER_38_492 ();
 sg13g2_decap_8 FILLER_38_529 ();
 sg13g2_decap_8 FILLER_38_536 ();
 sg13g2_decap_4 FILLER_38_543 ();
 sg13g2_decap_8 FILLER_38_558 ();
 sg13g2_decap_8 FILLER_38_565 ();
 sg13g2_fill_2 FILLER_38_572 ();
 sg13g2_decap_8 FILLER_38_600 ();
 sg13g2_fill_1 FILLER_38_607 ();
 sg13g2_fill_2 FILLER_38_612 ();
 sg13g2_fill_1 FILLER_38_631 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_decap_8 FILLER_38_669 ();
 sg13g2_decap_4 FILLER_38_676 ();
 sg13g2_fill_2 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_703 ();
 sg13g2_decap_8 FILLER_38_710 ();
 sg13g2_fill_2 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_719 ();
 sg13g2_fill_1 FILLER_38_747 ();
 sg13g2_fill_1 FILLER_38_752 ();
 sg13g2_fill_2 FILLER_38_762 ();
 sg13g2_fill_1 FILLER_38_764 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_4 FILLER_38_784 ();
 sg13g2_fill_2 FILLER_38_793 ();
 sg13g2_fill_1 FILLER_38_813 ();
 sg13g2_decap_4 FILLER_38_822 ();
 sg13g2_fill_1 FILLER_38_830 ();
 sg13g2_fill_1 FILLER_38_842 ();
 sg13g2_decap_4 FILLER_38_858 ();
 sg13g2_fill_2 FILLER_38_862 ();
 sg13g2_decap_8 FILLER_38_877 ();
 sg13g2_decap_8 FILLER_38_884 ();
 sg13g2_fill_2 FILLER_38_909 ();
 sg13g2_fill_1 FILLER_38_911 ();
 sg13g2_decap_8 FILLER_38_921 ();
 sg13g2_decap_8 FILLER_38_928 ();
 sg13g2_decap_8 FILLER_38_935 ();
 sg13g2_decap_8 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_949 ();
 sg13g2_decap_8 FILLER_38_956 ();
 sg13g2_decap_8 FILLER_38_963 ();
 sg13g2_decap_8 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_991 ();
 sg13g2_decap_8 FILLER_38_998 ();
 sg13g2_decap_8 FILLER_38_1005 ();
 sg13g2_decap_8 FILLER_38_1012 ();
 sg13g2_decap_4 FILLER_38_1019 ();
 sg13g2_fill_2 FILLER_38_1023 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_5 ();
 sg13g2_decap_4 FILLER_39_12 ();
 sg13g2_fill_2 FILLER_39_25 ();
 sg13g2_fill_1 FILLER_39_27 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_1 FILLER_39_211 ();
 sg13g2_fill_1 FILLER_39_230 ();
 sg13g2_fill_2 FILLER_39_308 ();
 sg13g2_fill_1 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_324 ();
 sg13g2_fill_2 FILLER_39_334 ();
 sg13g2_decap_8 FILLER_39_346 ();
 sg13g2_fill_2 FILLER_39_353 ();
 sg13g2_decap_4 FILLER_39_364 ();
 sg13g2_fill_2 FILLER_39_368 ();
 sg13g2_decap_4 FILLER_39_401 ();
 sg13g2_fill_2 FILLER_39_405 ();
 sg13g2_fill_2 FILLER_39_435 ();
 sg13g2_fill_1 FILLER_39_437 ();
 sg13g2_fill_1 FILLER_39_454 ();
 sg13g2_fill_2 FILLER_39_460 ();
 sg13g2_fill_1 FILLER_39_462 ();
 sg13g2_fill_2 FILLER_39_503 ();
 sg13g2_fill_1 FILLER_39_505 ();
 sg13g2_fill_2 FILLER_39_510 ();
 sg13g2_fill_1 FILLER_39_548 ();
 sg13g2_fill_1 FILLER_39_577 ();
 sg13g2_decap_8 FILLER_39_606 ();
 sg13g2_fill_1 FILLER_39_613 ();
 sg13g2_decap_4 FILLER_39_626 ();
 sg13g2_fill_2 FILLER_39_658 ();
 sg13g2_decap_4 FILLER_39_668 ();
 sg13g2_fill_1 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_fill_2 FILLER_39_735 ();
 sg13g2_fill_1 FILLER_39_737 ();
 sg13g2_fill_1 FILLER_39_762 ();
 sg13g2_fill_1 FILLER_39_787 ();
 sg13g2_fill_1 FILLER_39_802 ();
 sg13g2_fill_2 FILLER_39_808 ();
 sg13g2_fill_1 FILLER_39_818 ();
 sg13g2_decap_4 FILLER_39_824 ();
 sg13g2_fill_2 FILLER_39_852 ();
 sg13g2_fill_1 FILLER_39_854 ();
 sg13g2_fill_1 FILLER_39_860 ();
 sg13g2_fill_2 FILLER_39_866 ();
 sg13g2_decap_8 FILLER_39_896 ();
 sg13g2_decap_8 FILLER_39_903 ();
 sg13g2_decap_8 FILLER_39_910 ();
 sg13g2_decap_8 FILLER_39_917 ();
 sg13g2_decap_8 FILLER_39_924 ();
 sg13g2_decap_8 FILLER_39_931 ();
 sg13g2_decap_8 FILLER_39_938 ();
 sg13g2_decap_8 FILLER_39_945 ();
 sg13g2_decap_8 FILLER_39_952 ();
 sg13g2_decap_8 FILLER_39_959 ();
 sg13g2_decap_8 FILLER_39_966 ();
 sg13g2_decap_8 FILLER_39_973 ();
 sg13g2_decap_8 FILLER_39_980 ();
 sg13g2_decap_8 FILLER_39_987 ();
 sg13g2_decap_8 FILLER_39_994 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_8 FILLER_39_1008 ();
 sg13g2_decap_8 FILLER_39_1015 ();
 sg13g2_decap_8 FILLER_39_1022 ();
 sg13g2_decap_4 FILLER_40_4 ();
 sg13g2_fill_2 FILLER_40_8 ();
 sg13g2_fill_2 FILLER_40_42 ();
 sg13g2_fill_1 FILLER_40_44 ();
 sg13g2_fill_2 FILLER_40_85 ();
 sg13g2_fill_1 FILLER_40_87 ();
 sg13g2_decap_4 FILLER_40_92 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_fill_2 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_148 ();
 sg13g2_fill_2 FILLER_40_163 ();
 sg13g2_fill_2 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_348 ();
 sg13g2_decap_8 FILLER_40_355 ();
 sg13g2_decap_8 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_fill_1 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_380 ();
 sg13g2_fill_2 FILLER_40_390 ();
 sg13g2_fill_1 FILLER_40_392 ();
 sg13g2_fill_1 FILLER_40_402 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_40_423 ();
 sg13g2_decap_4 FILLER_40_430 ();
 sg13g2_fill_1 FILLER_40_434 ();
 sg13g2_fill_2 FILLER_40_439 ();
 sg13g2_fill_1 FILLER_40_441 ();
 sg13g2_decap_4 FILLER_40_474 ();
 sg13g2_decap_4 FILLER_40_483 ();
 sg13g2_fill_2 FILLER_40_487 ();
 sg13g2_decap_4 FILLER_40_498 ();
 sg13g2_fill_2 FILLER_40_524 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_fill_2 FILLER_40_560 ();
 sg13g2_fill_2 FILLER_40_584 ();
 sg13g2_fill_1 FILLER_40_586 ();
 sg13g2_fill_1 FILLER_40_603 ();
 sg13g2_decap_4 FILLER_40_607 ();
 sg13g2_fill_1 FILLER_40_611 ();
 sg13g2_fill_2 FILLER_40_624 ();
 sg13g2_decap_8 FILLER_40_632 ();
 sg13g2_decap_8 FILLER_40_639 ();
 sg13g2_decap_4 FILLER_40_646 ();
 sg13g2_fill_1 FILLER_40_650 ();
 sg13g2_fill_2 FILLER_40_655 ();
 sg13g2_decap_8 FILLER_40_699 ();
 sg13g2_decap_8 FILLER_40_706 ();
 sg13g2_decap_8 FILLER_40_713 ();
 sg13g2_decap_8 FILLER_40_720 ();
 sg13g2_decap_8 FILLER_40_727 ();
 sg13g2_decap_8 FILLER_40_734 ();
 sg13g2_fill_2 FILLER_40_741 ();
 sg13g2_fill_1 FILLER_40_743 ();
 sg13g2_fill_1 FILLER_40_749 ();
 sg13g2_fill_2 FILLER_40_756 ();
 sg13g2_decap_4 FILLER_40_777 ();
 sg13g2_fill_1 FILLER_40_781 ();
 sg13g2_decap_4 FILLER_40_826 ();
 sg13g2_fill_2 FILLER_40_848 ();
 sg13g2_fill_1 FILLER_40_850 ();
 sg13g2_fill_2 FILLER_40_868 ();
 sg13g2_decap_8 FILLER_40_879 ();
 sg13g2_decap_8 FILLER_40_886 ();
 sg13g2_decap_8 FILLER_40_893 ();
 sg13g2_decap_8 FILLER_40_900 ();
 sg13g2_decap_8 FILLER_40_907 ();
 sg13g2_decap_8 FILLER_40_914 ();
 sg13g2_decap_8 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_40_928 ();
 sg13g2_decap_8 FILLER_40_935 ();
 sg13g2_decap_8 FILLER_40_942 ();
 sg13g2_decap_8 FILLER_40_949 ();
 sg13g2_decap_8 FILLER_40_956 ();
 sg13g2_decap_8 FILLER_40_963 ();
 sg13g2_decap_8 FILLER_40_970 ();
 sg13g2_decap_8 FILLER_40_977 ();
 sg13g2_decap_8 FILLER_40_984 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_decap_8 FILLER_40_998 ();
 sg13g2_decap_8 FILLER_40_1005 ();
 sg13g2_decap_8 FILLER_40_1012 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_fill_2 FILLER_40_1026 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_fill_2 FILLER_41_36 ();
 sg13g2_fill_2 FILLER_41_47 ();
 sg13g2_fill_1 FILLER_41_49 ();
 sg13g2_fill_2 FILLER_41_55 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_fill_2 FILLER_41_133 ();
 sg13g2_fill_2 FILLER_41_139 ();
 sg13g2_fill_2 FILLER_41_160 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_fill_1 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_fill_1 FILLER_41_281 ();
 sg13g2_fill_2 FILLER_41_300 ();
 sg13g2_fill_1 FILLER_41_302 ();
 sg13g2_decap_4 FILLER_41_325 ();
 sg13g2_fill_2 FILLER_41_366 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_383 ();
 sg13g2_decap_4 FILLER_41_389 ();
 sg13g2_fill_2 FILLER_41_393 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_1 FILLER_41_435 ();
 sg13g2_decap_8 FILLER_41_487 ();
 sg13g2_decap_8 FILLER_41_494 ();
 sg13g2_decap_8 FILLER_41_501 ();
 sg13g2_decap_4 FILLER_41_508 ();
 sg13g2_decap_4 FILLER_41_539 ();
 sg13g2_fill_1 FILLER_41_570 ();
 sg13g2_fill_2 FILLER_41_598 ();
 sg13g2_decap_8 FILLER_41_622 ();
 sg13g2_decap_8 FILLER_41_629 ();
 sg13g2_decap_8 FILLER_41_636 ();
 sg13g2_fill_2 FILLER_41_643 ();
 sg13g2_fill_1 FILLER_41_653 ();
 sg13g2_decap_8 FILLER_41_660 ();
 sg13g2_decap_4 FILLER_41_667 ();
 sg13g2_decap_8 FILLER_41_675 ();
 sg13g2_decap_4 FILLER_41_682 ();
 sg13g2_decap_8 FILLER_41_712 ();
 sg13g2_fill_1 FILLER_41_766 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_818 ();
 sg13g2_decap_8 FILLER_41_825 ();
 sg13g2_fill_1 FILLER_41_832 ();
 sg13g2_fill_1 FILLER_41_841 ();
 sg13g2_fill_1 FILLER_41_849 ();
 sg13g2_decap_8 FILLER_41_891 ();
 sg13g2_decap_8 FILLER_41_898 ();
 sg13g2_decap_8 FILLER_41_905 ();
 sg13g2_decap_8 FILLER_41_912 ();
 sg13g2_decap_8 FILLER_41_919 ();
 sg13g2_decap_8 FILLER_41_926 ();
 sg13g2_decap_8 FILLER_41_933 ();
 sg13g2_decap_8 FILLER_41_940 ();
 sg13g2_decap_8 FILLER_41_947 ();
 sg13g2_decap_8 FILLER_41_954 ();
 sg13g2_decap_8 FILLER_41_961 ();
 sg13g2_decap_8 FILLER_41_968 ();
 sg13g2_decap_8 FILLER_41_975 ();
 sg13g2_decap_8 FILLER_41_982 ();
 sg13g2_decap_8 FILLER_41_989 ();
 sg13g2_decap_8 FILLER_41_996 ();
 sg13g2_decap_8 FILLER_41_1003 ();
 sg13g2_decap_8 FILLER_41_1010 ();
 sg13g2_decap_8 FILLER_41_1017 ();
 sg13g2_decap_4 FILLER_41_1024 ();
 sg13g2_fill_1 FILLER_41_1028 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_21 ();
 sg13g2_fill_1 FILLER_42_69 ();
 sg13g2_decap_4 FILLER_42_124 ();
 sg13g2_fill_2 FILLER_42_128 ();
 sg13g2_fill_2 FILLER_42_180 ();
 sg13g2_decap_8 FILLER_42_209 ();
 sg13g2_decap_4 FILLER_42_216 ();
 sg13g2_decap_8 FILLER_42_223 ();
 sg13g2_decap_8 FILLER_42_230 ();
 sg13g2_fill_2 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_decap_8 FILLER_42_244 ();
 sg13g2_fill_2 FILLER_42_251 ();
 sg13g2_fill_1 FILLER_42_253 ();
 sg13g2_decap_4 FILLER_42_299 ();
 sg13g2_decap_8 FILLER_42_312 ();
 sg13g2_decap_8 FILLER_42_319 ();
 sg13g2_fill_1 FILLER_42_348 ();
 sg13g2_decap_4 FILLER_42_363 ();
 sg13g2_fill_2 FILLER_42_405 ();
 sg13g2_fill_1 FILLER_42_407 ();
 sg13g2_fill_2 FILLER_42_445 ();
 sg13g2_fill_1 FILLER_42_447 ();
 sg13g2_fill_2 FILLER_42_476 ();
 sg13g2_fill_1 FILLER_42_478 ();
 sg13g2_decap_8 FILLER_42_506 ();
 sg13g2_fill_2 FILLER_42_513 ();
 sg13g2_fill_2 FILLER_42_533 ();
 sg13g2_decap_8 FILLER_42_544 ();
 sg13g2_decap_8 FILLER_42_551 ();
 sg13g2_decap_4 FILLER_42_585 ();
 sg13g2_fill_2 FILLER_42_589 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_fill_2 FILLER_42_798 ();
 sg13g2_fill_1 FILLER_42_800 ();
 sg13g2_fill_1 FILLER_42_828 ();
 sg13g2_fill_2 FILLER_42_875 ();
 sg13g2_decap_8 FILLER_42_886 ();
 sg13g2_decap_8 FILLER_42_893 ();
 sg13g2_decap_8 FILLER_42_900 ();
 sg13g2_decap_8 FILLER_42_907 ();
 sg13g2_decap_8 FILLER_42_914 ();
 sg13g2_decap_8 FILLER_42_921 ();
 sg13g2_decap_8 FILLER_42_928 ();
 sg13g2_decap_8 FILLER_42_935 ();
 sg13g2_decap_8 FILLER_42_942 ();
 sg13g2_decap_8 FILLER_42_949 ();
 sg13g2_decap_8 FILLER_42_956 ();
 sg13g2_decap_8 FILLER_42_963 ();
 sg13g2_decap_8 FILLER_42_970 ();
 sg13g2_decap_8 FILLER_42_977 ();
 sg13g2_decap_8 FILLER_42_984 ();
 sg13g2_decap_8 FILLER_42_991 ();
 sg13g2_decap_8 FILLER_42_998 ();
 sg13g2_decap_8 FILLER_42_1005 ();
 sg13g2_decap_8 FILLER_42_1012 ();
 sg13g2_decap_8 FILLER_42_1019 ();
 sg13g2_fill_2 FILLER_42_1026 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_2 FILLER_43_31 ();
 sg13g2_fill_1 FILLER_43_33 ();
 sg13g2_fill_2 FILLER_43_47 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_fill_1 FILLER_43_79 ();
 sg13g2_fill_1 FILLER_43_89 ();
 sg13g2_fill_2 FILLER_43_109 ();
 sg13g2_fill_1 FILLER_43_111 ();
 sg13g2_fill_1 FILLER_43_148 ();
 sg13g2_fill_1 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_decap_4 FILLER_43_205 ();
 sg13g2_fill_1 FILLER_43_246 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_fill_2 FILLER_43_298 ();
 sg13g2_decap_8 FILLER_43_316 ();
 sg13g2_decap_8 FILLER_43_323 ();
 sg13g2_fill_2 FILLER_43_351 ();
 sg13g2_fill_1 FILLER_43_353 ();
 sg13g2_decap_8 FILLER_43_359 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_fill_1 FILLER_43_392 ();
 sg13g2_fill_2 FILLER_43_417 ();
 sg13g2_fill_1 FILLER_43_419 ();
 sg13g2_decap_8 FILLER_43_438 ();
 sg13g2_fill_2 FILLER_43_445 ();
 sg13g2_fill_1 FILLER_43_456 ();
 sg13g2_decap_4 FILLER_43_482 ();
 sg13g2_fill_2 FILLER_43_486 ();
 sg13g2_decap_8 FILLER_43_563 ();
 sg13g2_decap_8 FILLER_43_570 ();
 sg13g2_fill_1 FILLER_43_577 ();
 sg13g2_decap_4 FILLER_43_587 ();
 sg13g2_fill_2 FILLER_43_591 ();
 sg13g2_fill_2 FILLER_43_604 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_fill_2 FILLER_43_622 ();
 sg13g2_fill_1 FILLER_43_624 ();
 sg13g2_decap_4 FILLER_43_638 ();
 sg13g2_decap_8 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_689 ();
 sg13g2_fill_2 FILLER_43_696 ();
 sg13g2_fill_1 FILLER_43_725 ();
 sg13g2_fill_1 FILLER_43_786 ();
 sg13g2_decap_8 FILLER_43_827 ();
 sg13g2_decap_8 FILLER_43_834 ();
 sg13g2_decap_8 FILLER_43_841 ();
 sg13g2_decap_8 FILLER_43_848 ();
 sg13g2_decap_8 FILLER_43_859 ();
 sg13g2_decap_8 FILLER_43_866 ();
 sg13g2_decap_8 FILLER_43_873 ();
 sg13g2_decap_8 FILLER_43_880 ();
 sg13g2_decap_8 FILLER_43_887 ();
 sg13g2_decap_8 FILLER_43_894 ();
 sg13g2_decap_8 FILLER_43_901 ();
 sg13g2_decap_8 FILLER_43_908 ();
 sg13g2_decap_8 FILLER_43_915 ();
 sg13g2_decap_8 FILLER_43_922 ();
 sg13g2_decap_8 FILLER_43_929 ();
 sg13g2_decap_8 FILLER_43_936 ();
 sg13g2_decap_8 FILLER_43_943 ();
 sg13g2_decap_8 FILLER_43_950 ();
 sg13g2_decap_8 FILLER_43_957 ();
 sg13g2_decap_8 FILLER_43_964 ();
 sg13g2_decap_8 FILLER_43_971 ();
 sg13g2_decap_8 FILLER_43_978 ();
 sg13g2_decap_8 FILLER_43_985 ();
 sg13g2_decap_8 FILLER_43_992 ();
 sg13g2_decap_8 FILLER_43_999 ();
 sg13g2_decap_8 FILLER_43_1006 ();
 sg13g2_decap_8 FILLER_43_1013 ();
 sg13g2_decap_8 FILLER_43_1020 ();
 sg13g2_fill_2 FILLER_43_1027 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_67 ();
 sg13g2_fill_1 FILLER_44_69 ();
 sg13g2_fill_1 FILLER_44_79 ();
 sg13g2_fill_2 FILLER_44_93 ();
 sg13g2_fill_1 FILLER_44_95 ();
 sg13g2_decap_4 FILLER_44_126 ();
 sg13g2_fill_1 FILLER_44_130 ();
 sg13g2_fill_2 FILLER_44_140 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_decap_4 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_207 ();
 sg13g2_fill_2 FILLER_44_217 ();
 sg13g2_fill_1 FILLER_44_228 ();
 sg13g2_fill_2 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_276 ();
 sg13g2_decap_4 FILLER_44_283 ();
 sg13g2_fill_2 FILLER_44_287 ();
 sg13g2_fill_1 FILLER_44_301 ();
 sg13g2_fill_2 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_347 ();
 sg13g2_decap_4 FILLER_44_357 ();
 sg13g2_fill_2 FILLER_44_361 ();
 sg13g2_decap_4 FILLER_44_369 ();
 sg13g2_fill_2 FILLER_44_373 ();
 sg13g2_decap_4 FILLER_44_381 ();
 sg13g2_fill_1 FILLER_44_385 ();
 sg13g2_fill_1 FILLER_44_423 ();
 sg13g2_decap_4 FILLER_44_434 ();
 sg13g2_fill_1 FILLER_44_477 ();
 sg13g2_decap_8 FILLER_44_493 ();
 sg13g2_fill_2 FILLER_44_500 ();
 sg13g2_fill_2 FILLER_44_529 ();
 sg13g2_fill_1 FILLER_44_558 ();
 sg13g2_fill_1 FILLER_44_586 ();
 sg13g2_fill_2 FILLER_44_605 ();
 sg13g2_fill_2 FILLER_44_625 ();
 sg13g2_decap_8 FILLER_44_652 ();
 sg13g2_fill_2 FILLER_44_715 ();
 sg13g2_fill_1 FILLER_44_717 ();
 sg13g2_fill_1 FILLER_44_722 ();
 sg13g2_fill_2 FILLER_44_732 ();
 sg13g2_decap_8 FILLER_44_737 ();
 sg13g2_fill_2 FILLER_44_744 ();
 sg13g2_decap_4 FILLER_44_749 ();
 sg13g2_fill_2 FILLER_44_780 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_4 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_815 ();
 sg13g2_decap_8 FILLER_44_822 ();
 sg13g2_decap_8 FILLER_44_829 ();
 sg13g2_decap_8 FILLER_44_836 ();
 sg13g2_decap_8 FILLER_44_843 ();
 sg13g2_decap_8 FILLER_44_850 ();
 sg13g2_decap_8 FILLER_44_857 ();
 sg13g2_decap_8 FILLER_44_864 ();
 sg13g2_decap_8 FILLER_44_871 ();
 sg13g2_decap_8 FILLER_44_878 ();
 sg13g2_decap_8 FILLER_44_885 ();
 sg13g2_decap_8 FILLER_44_892 ();
 sg13g2_decap_8 FILLER_44_899 ();
 sg13g2_decap_8 FILLER_44_906 ();
 sg13g2_decap_8 FILLER_44_913 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_decap_8 FILLER_44_927 ();
 sg13g2_decap_8 FILLER_44_934 ();
 sg13g2_decap_8 FILLER_44_941 ();
 sg13g2_decap_8 FILLER_44_948 ();
 sg13g2_decap_8 FILLER_44_955 ();
 sg13g2_decap_8 FILLER_44_962 ();
 sg13g2_decap_8 FILLER_44_969 ();
 sg13g2_decap_8 FILLER_44_976 ();
 sg13g2_decap_8 FILLER_44_983 ();
 sg13g2_decap_8 FILLER_44_990 ();
 sg13g2_decap_8 FILLER_44_997 ();
 sg13g2_decap_8 FILLER_44_1004 ();
 sg13g2_decap_8 FILLER_44_1011 ();
 sg13g2_decap_8 FILLER_44_1018 ();
 sg13g2_decap_4 FILLER_44_1025 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_11 ();
 sg13g2_fill_1 FILLER_45_22 ();
 sg13g2_fill_2 FILLER_45_32 ();
 sg13g2_fill_2 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_122 ();
 sg13g2_decap_8 FILLER_45_129 ();
 sg13g2_fill_2 FILLER_45_190 ();
 sg13g2_fill_2 FILLER_45_229 ();
 sg13g2_fill_1 FILLER_45_231 ();
 sg13g2_fill_1 FILLER_45_272 ();
 sg13g2_fill_2 FILLER_45_332 ();
 sg13g2_fill_1 FILLER_45_334 ();
 sg13g2_decap_4 FILLER_45_345 ();
 sg13g2_decap_8 FILLER_45_353 ();
 sg13g2_decap_4 FILLER_45_360 ();
 sg13g2_fill_1 FILLER_45_364 ();
 sg13g2_fill_2 FILLER_45_391 ();
 sg13g2_fill_1 FILLER_45_393 ();
 sg13g2_decap_4 FILLER_45_422 ();
 sg13g2_fill_2 FILLER_45_426 ();
 sg13g2_fill_2 FILLER_45_456 ();
 sg13g2_decap_4 FILLER_45_493 ();
 sg13g2_fill_2 FILLER_45_506 ();
 sg13g2_fill_1 FILLER_45_508 ();
 sg13g2_fill_2 FILLER_45_531 ();
 sg13g2_decap_8 FILLER_45_555 ();
 sg13g2_fill_1 FILLER_45_562 ();
 sg13g2_fill_2 FILLER_45_590 ();
 sg13g2_fill_1 FILLER_45_600 ();
 sg13g2_fill_2 FILLER_45_617 ();
 sg13g2_fill_1 FILLER_45_619 ();
 sg13g2_fill_2 FILLER_45_659 ();
 sg13g2_decap_8 FILLER_45_680 ();
 sg13g2_decap_8 FILLER_45_687 ();
 sg13g2_decap_8 FILLER_45_694 ();
 sg13g2_decap_8 FILLER_45_701 ();
 sg13g2_decap_8 FILLER_45_708 ();
 sg13g2_decap_8 FILLER_45_715 ();
 sg13g2_decap_8 FILLER_45_722 ();
 sg13g2_decap_8 FILLER_45_729 ();
 sg13g2_decap_8 FILLER_45_736 ();
 sg13g2_decap_8 FILLER_45_743 ();
 sg13g2_decap_8 FILLER_45_750 ();
 sg13g2_fill_2 FILLER_45_757 ();
 sg13g2_fill_1 FILLER_45_759 ();
 sg13g2_decap_8 FILLER_45_769 ();
 sg13g2_decap_8 FILLER_45_776 ();
 sg13g2_decap_8 FILLER_45_783 ();
 sg13g2_decap_8 FILLER_45_790 ();
 sg13g2_decap_8 FILLER_45_797 ();
 sg13g2_fill_1 FILLER_45_804 ();
 sg13g2_decap_8 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_821 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_8 FILLER_45_856 ();
 sg13g2_decap_8 FILLER_45_863 ();
 sg13g2_decap_8 FILLER_45_870 ();
 sg13g2_decap_8 FILLER_45_877 ();
 sg13g2_decap_8 FILLER_45_884 ();
 sg13g2_decap_8 FILLER_45_891 ();
 sg13g2_decap_8 FILLER_45_898 ();
 sg13g2_decap_8 FILLER_45_905 ();
 sg13g2_decap_8 FILLER_45_912 ();
 sg13g2_decap_8 FILLER_45_919 ();
 sg13g2_decap_8 FILLER_45_926 ();
 sg13g2_decap_8 FILLER_45_933 ();
 sg13g2_decap_8 FILLER_45_940 ();
 sg13g2_decap_8 FILLER_45_947 ();
 sg13g2_decap_8 FILLER_45_954 ();
 sg13g2_decap_8 FILLER_45_961 ();
 sg13g2_decap_8 FILLER_45_968 ();
 sg13g2_decap_8 FILLER_45_975 ();
 sg13g2_decap_8 FILLER_45_982 ();
 sg13g2_decap_8 FILLER_45_989 ();
 sg13g2_decap_8 FILLER_45_996 ();
 sg13g2_decap_8 FILLER_45_1003 ();
 sg13g2_decap_8 FILLER_45_1010 ();
 sg13g2_decap_8 FILLER_45_1017 ();
 sg13g2_decap_4 FILLER_45_1024 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_fill_1 FILLER_46_76 ();
 sg13g2_fill_2 FILLER_46_85 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_decap_4 FILLER_46_107 ();
 sg13g2_fill_1 FILLER_46_111 ();
 sg13g2_decap_8 FILLER_46_121 ();
 sg13g2_fill_2 FILLER_46_128 ();
 sg13g2_fill_1 FILLER_46_165 ();
 sg13g2_fill_2 FILLER_46_211 ();
 sg13g2_decap_8 FILLER_46_235 ();
 sg13g2_decap_8 FILLER_46_242 ();
 sg13g2_fill_1 FILLER_46_249 ();
 sg13g2_fill_2 FILLER_46_278 ();
 sg13g2_fill_2 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_46_358 ();
 sg13g2_fill_1 FILLER_46_360 ();
 sg13g2_decap_8 FILLER_46_380 ();
 sg13g2_decap_8 FILLER_46_387 ();
 sg13g2_decap_4 FILLER_46_394 ();
 sg13g2_fill_2 FILLER_46_398 ();
 sg13g2_fill_1 FILLER_46_413 ();
 sg13g2_fill_2 FILLER_46_424 ();
 sg13g2_fill_1 FILLER_46_426 ();
 sg13g2_decap_4 FILLER_46_436 ();
 sg13g2_fill_2 FILLER_46_449 ();
 sg13g2_fill_1 FILLER_46_451 ();
 sg13g2_decap_4 FILLER_46_462 ();
 sg13g2_fill_2 FILLER_46_466 ();
 sg13g2_fill_2 FILLER_46_542 ();
 sg13g2_fill_1 FILLER_46_571 ();
 sg13g2_fill_1 FILLER_46_590 ();
 sg13g2_fill_2 FILLER_46_633 ();
 sg13g2_fill_1 FILLER_46_657 ();
 sg13g2_decap_8 FILLER_46_682 ();
 sg13g2_fill_1 FILLER_46_689 ();
 sg13g2_decap_4 FILLER_46_694 ();
 sg13g2_fill_2 FILLER_46_698 ();
 sg13g2_decap_8 FILLER_46_704 ();
 sg13g2_decap_8 FILLER_46_711 ();
 sg13g2_decap_8 FILLER_46_718 ();
 sg13g2_decap_8 FILLER_46_725 ();
 sg13g2_decap_8 FILLER_46_732 ();
 sg13g2_decap_8 FILLER_46_739 ();
 sg13g2_decap_8 FILLER_46_746 ();
 sg13g2_decap_8 FILLER_46_753 ();
 sg13g2_decap_8 FILLER_46_760 ();
 sg13g2_decap_8 FILLER_46_767 ();
 sg13g2_decap_8 FILLER_46_774 ();
 sg13g2_decap_8 FILLER_46_781 ();
 sg13g2_decap_8 FILLER_46_788 ();
 sg13g2_decap_8 FILLER_46_795 ();
 sg13g2_decap_8 FILLER_46_802 ();
 sg13g2_decap_8 FILLER_46_809 ();
 sg13g2_decap_8 FILLER_46_816 ();
 sg13g2_decap_8 FILLER_46_823 ();
 sg13g2_decap_8 FILLER_46_830 ();
 sg13g2_decap_8 FILLER_46_837 ();
 sg13g2_decap_8 FILLER_46_844 ();
 sg13g2_decap_8 FILLER_46_851 ();
 sg13g2_decap_8 FILLER_46_858 ();
 sg13g2_decap_8 FILLER_46_865 ();
 sg13g2_decap_8 FILLER_46_872 ();
 sg13g2_decap_8 FILLER_46_879 ();
 sg13g2_decap_8 FILLER_46_886 ();
 sg13g2_decap_8 FILLER_46_893 ();
 sg13g2_decap_8 FILLER_46_900 ();
 sg13g2_decap_8 FILLER_46_907 ();
 sg13g2_decap_8 FILLER_46_914 ();
 sg13g2_decap_8 FILLER_46_921 ();
 sg13g2_decap_8 FILLER_46_928 ();
 sg13g2_decap_8 FILLER_46_935 ();
 sg13g2_decap_8 FILLER_46_942 ();
 sg13g2_decap_8 FILLER_46_949 ();
 sg13g2_decap_8 FILLER_46_956 ();
 sg13g2_decap_8 FILLER_46_963 ();
 sg13g2_decap_8 FILLER_46_970 ();
 sg13g2_decap_8 FILLER_46_977 ();
 sg13g2_decap_8 FILLER_46_984 ();
 sg13g2_decap_8 FILLER_46_991 ();
 sg13g2_decap_8 FILLER_46_998 ();
 sg13g2_decap_8 FILLER_46_1005 ();
 sg13g2_decap_8 FILLER_46_1012 ();
 sg13g2_decap_8 FILLER_46_1019 ();
 sg13g2_fill_2 FILLER_46_1026 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_17 ();
 sg13g2_decap_4 FILLER_47_24 ();
 sg13g2_fill_2 FILLER_47_28 ();
 sg13g2_fill_2 FILLER_47_47 ();
 sg13g2_fill_1 FILLER_47_90 ();
 sg13g2_fill_2 FILLER_47_119 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_decap_4 FILLER_47_212 ();
 sg13g2_decap_8 FILLER_47_221 ();
 sg13g2_decap_4 FILLER_47_228 ();
 sg13g2_fill_1 FILLER_47_232 ();
 sg13g2_decap_4 FILLER_47_246 ();
 sg13g2_fill_2 FILLER_47_250 ();
 sg13g2_fill_2 FILLER_47_266 ();
 sg13g2_decap_4 FILLER_47_285 ();
 sg13g2_fill_1 FILLER_47_289 ();
 sg13g2_fill_2 FILLER_47_322 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_fill_2 FILLER_47_431 ();
 sg13g2_fill_2 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_480 ();
 sg13g2_decap_8 FILLER_47_487 ();
 sg13g2_decap_8 FILLER_47_494 ();
 sg13g2_decap_8 FILLER_47_501 ();
 sg13g2_decap_8 FILLER_47_508 ();
 sg13g2_decap_8 FILLER_47_515 ();
 sg13g2_fill_2 FILLER_47_522 ();
 sg13g2_fill_1 FILLER_47_524 ();
 sg13g2_fill_2 FILLER_47_529 ();
 sg13g2_decap_8 FILLER_47_536 ();
 sg13g2_decap_8 FILLER_47_543 ();
 sg13g2_decap_8 FILLER_47_550 ();
 sg13g2_decap_8 FILLER_47_557 ();
 sg13g2_decap_4 FILLER_47_564 ();
 sg13g2_decap_4 FILLER_47_585 ();
 sg13g2_fill_1 FILLER_47_589 ();
 sg13g2_fill_2 FILLER_47_596 ();
 sg13g2_fill_2 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_709 ();
 sg13g2_decap_8 FILLER_47_716 ();
 sg13g2_decap_8 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_730 ();
 sg13g2_decap_8 FILLER_47_737 ();
 sg13g2_decap_8 FILLER_47_744 ();
 sg13g2_decap_8 FILLER_47_751 ();
 sg13g2_decap_8 FILLER_47_758 ();
 sg13g2_decap_8 FILLER_47_765 ();
 sg13g2_decap_8 FILLER_47_772 ();
 sg13g2_decap_8 FILLER_47_779 ();
 sg13g2_decap_8 FILLER_47_786 ();
 sg13g2_decap_8 FILLER_47_793 ();
 sg13g2_decap_8 FILLER_47_800 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_decap_8 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_821 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_835 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_decap_8 FILLER_47_856 ();
 sg13g2_decap_8 FILLER_47_863 ();
 sg13g2_decap_8 FILLER_47_870 ();
 sg13g2_decap_8 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_47_884 ();
 sg13g2_decap_8 FILLER_47_891 ();
 sg13g2_decap_8 FILLER_47_898 ();
 sg13g2_decap_8 FILLER_47_905 ();
 sg13g2_decap_8 FILLER_47_912 ();
 sg13g2_decap_8 FILLER_47_919 ();
 sg13g2_decap_8 FILLER_47_926 ();
 sg13g2_decap_8 FILLER_47_933 ();
 sg13g2_decap_8 FILLER_47_940 ();
 sg13g2_decap_8 FILLER_47_947 ();
 sg13g2_decap_8 FILLER_47_954 ();
 sg13g2_decap_8 FILLER_47_961 ();
 sg13g2_decap_8 FILLER_47_968 ();
 sg13g2_decap_8 FILLER_47_975 ();
 sg13g2_decap_8 FILLER_47_982 ();
 sg13g2_decap_8 FILLER_47_989 ();
 sg13g2_decap_8 FILLER_47_996 ();
 sg13g2_decap_8 FILLER_47_1003 ();
 sg13g2_decap_8 FILLER_47_1010 ();
 sg13g2_decap_8 FILLER_47_1017 ();
 sg13g2_fill_1 FILLER_47_1024 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_fill_2 FILLER_48_35 ();
 sg13g2_fill_1 FILLER_48_37 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_fill_1 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_178 ();
 sg13g2_fill_2 FILLER_48_276 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_1 FILLER_48_338 ();
 sg13g2_fill_2 FILLER_48_449 ();
 sg13g2_decap_8 FILLER_48_488 ();
 sg13g2_decap_8 FILLER_48_495 ();
 sg13g2_decap_8 FILLER_48_502 ();
 sg13g2_decap_8 FILLER_48_509 ();
 sg13g2_decap_8 FILLER_48_516 ();
 sg13g2_decap_8 FILLER_48_523 ();
 sg13g2_decap_8 FILLER_48_530 ();
 sg13g2_decap_8 FILLER_48_537 ();
 sg13g2_decap_8 FILLER_48_544 ();
 sg13g2_decap_8 FILLER_48_551 ();
 sg13g2_decap_8 FILLER_48_558 ();
 sg13g2_decap_4 FILLER_48_565 ();
 sg13g2_fill_2 FILLER_48_569 ();
 sg13g2_fill_2 FILLER_48_625 ();
 sg13g2_fill_1 FILLER_48_627 ();
 sg13g2_decap_8 FILLER_48_655 ();
 sg13g2_decap_4 FILLER_48_662 ();
 sg13g2_fill_2 FILLER_48_666 ();
 sg13g2_fill_2 FILLER_48_695 ();
 sg13g2_fill_1 FILLER_48_697 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_48_931 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_945 ();
 sg13g2_decap_8 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_959 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_4 FILLER_49_53 ();
 sg13g2_fill_2 FILLER_49_57 ();
 sg13g2_decap_4 FILLER_49_64 ();
 sg13g2_fill_2 FILLER_49_68 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_fill_2 FILLER_49_142 ();
 sg13g2_fill_2 FILLER_49_170 ();
 sg13g2_fill_1 FILLER_49_172 ();
 sg13g2_decap_4 FILLER_49_192 ();
 sg13g2_decap_4 FILLER_49_214 ();
 sg13g2_fill_1 FILLER_49_218 ();
 sg13g2_fill_2 FILLER_49_238 ();
 sg13g2_fill_1 FILLER_49_240 ();
 sg13g2_decap_8 FILLER_49_250 ();
 sg13g2_decap_8 FILLER_49_257 ();
 sg13g2_decap_4 FILLER_49_264 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_fill_1 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_313 ();
 sg13g2_decap_4 FILLER_49_320 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_fill_2 FILLER_49_340 ();
 sg13g2_fill_1 FILLER_49_351 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_fill_2 FILLER_49_382 ();
 sg13g2_fill_1 FILLER_49_384 ();
 sg13g2_fill_2 FILLER_49_412 ();
 sg13g2_fill_1 FILLER_49_423 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_4 FILLER_49_452 ();
 sg13g2_fill_1 FILLER_49_456 ();
 sg13g2_decap_8 FILLER_49_470 ();
 sg13g2_decap_8 FILLER_49_477 ();
 sg13g2_decap_8 FILLER_49_484 ();
 sg13g2_decap_8 FILLER_49_491 ();
 sg13g2_decap_8 FILLER_49_498 ();
 sg13g2_decap_8 FILLER_49_505 ();
 sg13g2_decap_8 FILLER_49_512 ();
 sg13g2_decap_8 FILLER_49_519 ();
 sg13g2_decap_8 FILLER_49_526 ();
 sg13g2_decap_8 FILLER_49_533 ();
 sg13g2_decap_8 FILLER_49_540 ();
 sg13g2_decap_8 FILLER_49_547 ();
 sg13g2_decap_8 FILLER_49_554 ();
 sg13g2_decap_8 FILLER_49_561 ();
 sg13g2_fill_2 FILLER_49_568 ();
 sg13g2_fill_1 FILLER_49_570 ();
 sg13g2_decap_8 FILLER_49_584 ();
 sg13g2_decap_8 FILLER_49_591 ();
 sg13g2_decap_4 FILLER_49_598 ();
 sg13g2_decap_4 FILLER_49_608 ();
 sg13g2_fill_2 FILLER_49_612 ();
 sg13g2_decap_4 FILLER_49_632 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_decap_8 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_662 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_decap_8 FILLER_49_683 ();
 sg13g2_decap_8 FILLER_49_690 ();
 sg13g2_decap_8 FILLER_49_697 ();
 sg13g2_decap_8 FILLER_49_704 ();
 sg13g2_decap_8 FILLER_49_711 ();
 sg13g2_decap_8 FILLER_49_718 ();
 sg13g2_decap_8 FILLER_49_725 ();
 sg13g2_decap_8 FILLER_49_732 ();
 sg13g2_decap_8 FILLER_49_739 ();
 sg13g2_decap_8 FILLER_49_746 ();
 sg13g2_decap_8 FILLER_49_753 ();
 sg13g2_decap_8 FILLER_49_760 ();
 sg13g2_decap_8 FILLER_49_767 ();
 sg13g2_decap_8 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_781 ();
 sg13g2_decap_8 FILLER_49_788 ();
 sg13g2_decap_8 FILLER_49_795 ();
 sg13g2_decap_8 FILLER_49_802 ();
 sg13g2_decap_8 FILLER_49_809 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_decap_8 FILLER_49_823 ();
 sg13g2_decap_8 FILLER_49_830 ();
 sg13g2_decap_8 FILLER_49_837 ();
 sg13g2_decap_8 FILLER_49_844 ();
 sg13g2_decap_8 FILLER_49_851 ();
 sg13g2_decap_8 FILLER_49_858 ();
 sg13g2_decap_8 FILLER_49_865 ();
 sg13g2_decap_8 FILLER_49_872 ();
 sg13g2_decap_8 FILLER_49_879 ();
 sg13g2_decap_8 FILLER_49_886 ();
 sg13g2_decap_8 FILLER_49_893 ();
 sg13g2_decap_8 FILLER_49_900 ();
 sg13g2_decap_8 FILLER_49_907 ();
 sg13g2_decap_8 FILLER_49_914 ();
 sg13g2_decap_8 FILLER_49_921 ();
 sg13g2_decap_8 FILLER_49_928 ();
 sg13g2_decap_8 FILLER_49_935 ();
 sg13g2_decap_8 FILLER_49_942 ();
 sg13g2_decap_8 FILLER_49_949 ();
 sg13g2_decap_8 FILLER_49_956 ();
 sg13g2_decap_8 FILLER_49_963 ();
 sg13g2_decap_8 FILLER_49_970 ();
 sg13g2_decap_8 FILLER_49_977 ();
 sg13g2_decap_8 FILLER_49_984 ();
 sg13g2_decap_8 FILLER_49_991 ();
 sg13g2_decap_8 FILLER_49_998 ();
 sg13g2_decap_8 FILLER_49_1005 ();
 sg13g2_decap_8 FILLER_49_1012 ();
 sg13g2_decap_8 FILLER_49_1019 ();
 sg13g2_fill_2 FILLER_49_1026 ();
 sg13g2_fill_1 FILLER_49_1028 ();
 assign uio_out[7] = net41;
endmodule
