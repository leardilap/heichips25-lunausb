* NGSPICE file created from heichips25_usb_cdc.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

.subckt heichips25_usb_cdc VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] usb_dn_en_o usb_dn_rx_i usb_dn_tx_o usb_dp_en_o usb_dp_rx_i
+ usb_dp_tx_o
XFILLER_39_211 VPWR VGND sg13g2_fill_1
X_3155_ _1235_ net100 _1230_ VPWR VGND sg13g2_nand2_1
XFILLER_28_929 VPWR VGND sg13g2_fill_1
X_3086_ _1198_ net240 net606 VPWR VGND sg13g2_nand2_1
X_2106_ VPWR _1984_ net382 VGND sg13g2_inv_1
XFILLER_36_940 VPWR VGND sg13g2_decap_8
X_2037_ VPWR _1916_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[1\] VGND sg13g2_inv_1
XFILLER_22_155 VPWR VGND sg13g2_fill_1
X_3988_ net931 _1999_ _2003_ _0954_ _1872_ VPWR VGND sg13g2_nor4_1
X_2939_ _1117_ net87 _1110_ VPWR VGND sg13g2_nand2_1
Xhold362 net29 VPWR VGND net404 sg13g2_dlygate4sd3_1
XFILLER_2_516 VPWR VGND sg13g2_decap_8
Xhold351 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[9\] VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold340 _0053_ VPWR VGND net382 sg13g2_dlygate4sd3_1
Xhold384 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[26\] VPWR VGND
+ net426 sg13g2_dlygate4sd3_1
Xhold373 _0055_ VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold395 _0115_ VPWR VGND net437 sg13g2_dlygate4sd3_1
Xfanout842 net1029 net842 VPWR VGND sg13g2_buf_8
Xfanout820 net821 net820 VPWR VGND sg13g2_buf_8
Xfanout831 u_usb_cdc.u_sie.phy_state_q\[10\] net831 VPWR VGND sg13g2_buf_8
XFILLER_46_704 VPWR VGND sg13g2_decap_8
XFILLER_19_929 VPWR VGND sg13g2_fill_1
XFILLER_42_921 VPWR VGND sg13g2_decap_8
XFILLER_42_998 VPWR VGND sg13g2_decap_8
XFILLER_6_800 VPWR VGND sg13g2_decap_8
XFILLER_6_877 VPWR VGND sg13g2_decap_8
XFILLER_1_582 VPWR VGND sg13g2_decap_8
XFILLER_3_1018 VPWR VGND sg13g2_decap_8
XFILLER_37_715 VPWR VGND sg13g2_fill_1
XFILLER_18_951 VPWR VGND sg13g2_decap_8
X_3911_ _1805_ net829 _2003_ VPWR VGND sg13g2_nand2_1
XFILLER_33_965 VPWR VGND sg13g2_decap_8
X_3842_ _1764_ VPWR _0390_ VGND _1765_ _1766_ sg13g2_o21ai_1
XFILLER_20_604 VPWR VGND sg13g2_fill_2
XFILLER_20_626 VPWR VGND sg13g2_fill_1
XFILLER_20_637 VPWR VGND sg13g2_fill_2
XFILLER_32_497 VPWR VGND sg13g2_decap_8
X_3773_ net291 _1716_ _1717_ VPWR VGND sg13g2_nor2_1
X_2724_ VGND VPWR _1893_ net38 _1975_ net829 sg13g2_a21oi_2
X_2655_ _0924_ _0925_ _0923_ _0029_ VPWR VGND sg13g2_nand3_1
X_4325_ net687 VGND VPWR _0327_ u_usb_cdc.u_sie.crc16_q\[4\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_2586_ _0868_ net840 net595 VPWR VGND sg13g2_nand2_1
X_4256_ net643 VGND VPWR _0258_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[3\]
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_41_1024 VPWR VGND sg13g2_decap_4
X_3207_ net809 net807 _1279_ VPWR VGND sg13g2_nor2_2
X_4187_ net646 VGND VPWR net315 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[23\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3138_ _1225_ VPWR _0227_ VGND _1899_ net627 sg13g2_o21ai_1
X_3069_ _1189_ net176 net609 VPWR VGND sg13g2_nand2_1
XFILLER_42_239 VPWR VGND sg13g2_fill_1
XFILLER_24_954 VPWR VGND sg13g2_fill_2
XFILLER_10_125 VPWR VGND sg13g2_decap_8
XFILLER_3_836 VPWR VGND sg13g2_decap_8
XFILLER_2_302 VPWR VGND sg13g2_fill_2
Xhold170 _0423_ VPWR VGND net212 sg13g2_dlygate4sd3_1
XFILLER_5_4 VPWR VGND sg13g2_fill_2
XFILLER_2_357 VPWR VGND sg13g2_decap_8
Xhold181 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[56\] VPWR
+ VGND net223 sg13g2_dlygate4sd3_1
Xhold192 u_usb_cdc.dp_pu_o VPWR VGND net234 sg13g2_dlygate4sd3_1
Xfanout650 net652 net650 VPWR VGND sg13g2_buf_8
Xfanout661 net664 net661 VPWR VGND sg13g2_buf_8
Xfanout694 net697 net694 VPWR VGND sg13g2_buf_8
Xfanout672 net675 net672 VPWR VGND sg13g2_buf_8
Xfanout683 net685 net683 VPWR VGND sg13g2_buf_8
XFILLER_19_759 VPWR VGND sg13g2_fill_1
XFILLER_34_729 VPWR VGND sg13g2_fill_2
XFILLER_15_998 VPWR VGND sg13g2_decap_8
X_2440_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[1\] _0547_ _0738_ VPWR VGND sg13g2_nor2_1
X_2371_ _0550_ _0670_ _0671_ VPWR VGND sg13g2_nor2_1
XFILLER_38_4 VPWR VGND sg13g2_fill_1
X_4110_ net669 VGND VPWR net457 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[30\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_25_1019 VPWR VGND sg13g2_decap_8
X_4041_ net678 VGND VPWR net867 u_usb_cdc.u_ctrl_endp.state_q\[5\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_37_578 VPWR VGND sg13g2_decap_8
XFILLER_37_589 VPWR VGND sg13g2_fill_2
XFILLER_33_795 VPWR VGND sg13g2_decap_4
X_3825_ _1738_ _1753_ _1754_ VPWR VGND sg13g2_nor2_1
XFILLER_20_434 VPWR VGND sg13g2_decap_8
XFILLER_20_478 VPWR VGND sg13g2_decap_8
X_3756_ _0889_ _1692_ net1011 _1702_ VPWR VGND sg13g2_nand3_1
X_2707_ _0962_ _0964_ _0961_ _0965_ VPWR VGND sg13g2_nand3_1
X_3687_ net790 VPWR _1657_ VGND _1655_ _1656_ sg13g2_o21ai_1
X_2638_ _0910_ net592 _0909_ net595 net975 VPWR VGND sg13g2_a22oi_1
X_2569_ _0626_ _0628_ _0856_ VPWR VGND sg13g2_nor2_1
X_4308_ net691 VGND VPWR net238 u_usb_cdc.u_sie.addr_q\[4\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_4239_ net642 VGND VPWR _0242_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\]
+ clknet_leaf_4_clk sg13g2_dfrbpq_2
XFILLER_16_707 VPWR VGND sg13g2_fill_2
XFILLER_28_567 VPWR VGND sg13g2_fill_1
XFILLER_15_206 VPWR VGND sg13g2_decap_8
XFILLER_8_917 VPWR VGND sg13g2_decap_8
XFILLER_12_979 VPWR VGND sg13g2_decap_8
XFILLER_48_1008 VPWR VGND sg13g2_decap_8
XFILLER_3_633 VPWR VGND sg13g2_decap_8
XFILLER_47_821 VPWR VGND sg13g2_decap_8
XFILLER_19_512 VPWR VGND sg13g2_fill_2
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_47_898 VPWR VGND sg13g2_decap_8
XFILLER_34_559 VPWR VGND sg13g2_fill_2
XFILLER_14_250 VPWR VGND sg13g2_decap_8
XFILLER_14_261 VPWR VGND sg13g2_fill_2
XFILLER_15_795 VPWR VGND sg13g2_fill_2
XFILLER_9_77 VPWR VGND sg13g2_fill_1
X_3610_ _1583_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[67\] net626
+ VPWR VGND sg13g2_nand2_1
X_3541_ VPWR _1517_ _1516_ VGND sg13g2_inv_1
XFILLER_7_983 VPWR VGND sg13g2_decap_8
XFILLER_6_471 VPWR VGND sg13g2_decap_8
X_3472_ VGND VPWR u_usb_cdc.u_sie.delay_cnt_q\[0\] net742 _1470_ net507 sg13g2_a21oi_1
XFILLER_43_2 VPWR VGND sg13g2_fill_1
X_2423_ _0699_ _0714_ _0721_ VPWR VGND sg13g2_nor2_1
X_2354_ VGND VPWR _0654_ _0649_ net779 sg13g2_or2_1
X_2285_ _0587_ _1997_ _0586_ VPWR VGND sg13g2_nand2b_1
X_4024_ net676 VGND VPWR net972 u_usb_cdc.u_ctrl_endp.req_q\[4\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_2
X_3808_ VGND VPWR net740 net318 _0381_ _1741_ sg13g2_a21oi_1
X_3739_ net751 net843 _0602_ _0362_ VPWR VGND sg13g2_mux2_1
XFILLER_0_647 VPWR VGND sg13g2_decap_8
XFILLER_28_331 VPWR VGND sg13g2_fill_1
XFILLER_44_857 VPWR VGND sg13g2_decap_8
XFILLER_43_323 VPWR VGND sg13g2_decap_8
XFILLER_28_397 VPWR VGND sg13g2_fill_1
XFILLER_31_507 VPWR VGND sg13g2_decap_8
XFILLER_24_570 VPWR VGND sg13g2_fill_1
XFILLER_12_754 VPWR VGND sg13g2_fill_2
XFILLER_34_96 VPWR VGND sg13g2_fill_1
XFILLER_8_769 VPWR VGND sg13g2_decap_8
XFILLER_4_942 VPWR VGND sg13g2_decap_8
XFILLER_3_452 VPWR VGND sg13g2_decap_8
XFILLER_3_441 VPWR VGND sg13g2_fill_2
XFILLER_38_128 VPWR VGND sg13g2_decap_8
X_2070_ VPWR _1949_ net502 VGND sg13g2_inv_1
XFILLER_38_139 VPWR VGND sg13g2_fill_1
XFILLER_19_375 VPWR VGND sg13g2_fill_2
XFILLER_19_397 VPWR VGND sg13g2_fill_2
XFILLER_35_835 VPWR VGND sg13g2_fill_1
X_2972_ _1041_ net997 _1055_ _0159_ VPWR VGND sg13g2_mux2_1
Xhold703 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ VPWR VGND net1021 sg13g2_dlygate4sd3_1
Xhold736 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[0\] VPWR
+ VGND net1054 sg13g2_dlygate4sd3_1
Xhold725 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[1\] VPWR VGND net1043 sg13g2_dlygate4sd3_1
Xhold714 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ VPWR VGND net1032 sg13g2_dlygate4sd3_1
X_3524_ _1500_ _1494_ _1499_ net626 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[64\]
+ VPWR VGND sg13g2_a22oi_1
Xhold747 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\] VPWR VGND
+ net1065 sg13g2_dlygate4sd3_1
X_3455_ u_usb_cdc.u_ctrl_endp.addr_dd\[2\] u_usb_cdc.u_ctrl_endp.addr_dd\[5\] u_usb_cdc.u_ctrl_endp.addr_dd\[4\]
+ u_usb_cdc.u_ctrl_endp.addr_dd\[6\] _1457_ VPWR VGND sg13g2_nor4_1
X_2406_ net784 _0654_ _0661_ _0704_ _0706_ VPWR VGND sg13g2_nor4_1
X_3386_ VGND VPWR net567 _1411_ _0289_ _1410_ sg13g2_a21oi_1
X_2337_ net588 _0637_ _0638_ VPWR VGND sg13g2_nor2_2
X_2268_ net706 VPWR _0570_ VGND _0568_ _0569_ sg13g2_o21ai_1
XFILLER_26_824 VPWR VGND sg13g2_decap_8
X_4007_ _1886_ net85 _1885_ VPWR VGND sg13g2_nand2_1
X_2199_ u_usb_cdc.u_sie.data_q\[6\] net540 _0501_ VPWR VGND sg13g2_xor2_1
XFILLER_41_849 VPWR VGND sg13g2_fill_1
XFILLER_40_348 VPWR VGND sg13g2_decap_8
XFILLER_0_444 VPWR VGND sg13g2_decap_8
XFILLER_1_967 VPWR VGND sg13g2_decap_8
XFILLER_49_949 VPWR VGND sg13g2_decap_8
Xhold30 _0129_ VPWR VGND net72 sg13g2_dlygate4sd3_1
Xhold41 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[40\] VPWR VGND
+ net83 sg13g2_dlygate4sd3_1
Xhold52 _0104_ VPWR VGND net94 sg13g2_dlygate4sd3_1
Xhold63 _0175_ VPWR VGND net105 sg13g2_dlygate4sd3_1
Xhold74 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[70\] VPWR VGND
+ net116 sg13g2_dlygate4sd3_1
XFILLER_29_640 VPWR VGND sg13g2_fill_1
Xhold96 _0094_ VPWR VGND net138 sg13g2_dlygate4sd3_1
Xhold85 _0135_ VPWR VGND net127 sg13g2_dlygate4sd3_1
XFILLER_17_857 VPWR VGND sg13g2_fill_1
XFILLER_28_161 VPWR VGND sg13g2_decap_8
XFILLER_16_334 VPWR VGND sg13g2_decap_8
XFILLER_12_540 VPWR VGND sg13g2_decap_4
XFILLER_40_893 VPWR VGND sg13g2_decap_8
XFILLER_8_533 VPWR VGND sg13g2_fill_1
XFILLER_6_45 VPWR VGND sg13g2_decap_4
X_3240_ VGND VPWR _1309_ net63 net812 sg13g2_or2_1
XFILLER_3_293 VPWR VGND sg13g2_decap_8
X_3171_ _1244_ _1246_ _1243_ _1247_ VPWR VGND sg13g2_nand3_1
X_2122_ _2000_ _1993_ net623 VPWR VGND sg13g2_nand2_1
XFILLER_39_437 VPWR VGND sg13g2_fill_1
X_2053_ _1932_ net842 VPWR VGND sg13g2_inv_2
XFILLER_23_805 VPWR VGND sg13g2_fill_2
XFILLER_34_120 VPWR VGND sg13g2_fill_2
XFILLER_22_315 VPWR VGND sg13g2_decap_8
X_2955_ net430 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ _1121_ _0148_ VPWR VGND sg13g2_mux2_1
X_2886_ _1094_ VPWR _0105_ VGND net824 _1095_ sg13g2_o21ai_1
Xhold511 _0001_ VPWR VGND net553 sg13g2_dlygate4sd3_1
Xhold500 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q
+ VPWR VGND net542 sg13g2_dlygate4sd3_1
X_3507_ _0336_ net572 _1950_ net575 _1940_ VPWR VGND sg13g2_a22oi_1
Xhold533 _0068_ VPWR VGND net851 sg13g2_dlygate4sd3_1
Xhold544 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[6\] VPWR VGND net862 sg13g2_dlygate4sd3_1
Xhold522 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq
+ VPWR VGND net564 sg13g2_dlygate4sd3_1
Xhold566 u_usb_cdc.u_ctrl_endp.class_q VPWR VGND net884 sg13g2_dlygate4sd3_1
Xhold577 _0244_ VPWR VGND net895 sg13g2_dlygate4sd3_1
Xhold555 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[7\] VPWR VGND net873 sg13g2_dlygate4sd3_1
Xhold588 u_usb_cdc.u_ctrl_endp.req_q\[6\] VPWR VGND net906 sg13g2_dlygate4sd3_1
XFILLER_44_1011 VPWR VGND sg13g2_decap_8
Xhold599 _0291_ VPWR VGND net917 sg13g2_dlygate4sd3_1
X_3438_ net764 net1002 net582 _0305_ VPWR VGND sg13g2_mux2_1
X_3369_ net920 _1399_ _1400_ VPWR VGND sg13g2_nor2_1
XFILLER_38_492 VPWR VGND sg13g2_fill_2
XFILLER_14_827 VPWR VGND sg13g2_decap_4
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_5_514 VPWR VGND sg13g2_fill_2
XFILLER_31_20 VPWR VGND sg13g2_fill_2
XFILLER_31_31 VPWR VGND sg13g2_decap_4
Xoutput31 net31 uo_out[2] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uio_oe[6] VPWR VGND sg13g2_buf_1
XFILLER_0_263 VPWR VGND sg13g2_fill_2
XFILLER_1_764 VPWR VGND sg13g2_decap_8
XFILLER_49_746 VPWR VGND sg13g2_decap_8
XFILLER_48_278 VPWR VGND sg13g2_fill_1
XFILLER_45_996 VPWR VGND sg13g2_decap_8
XFILLER_17_676 VPWR VGND sg13g2_fill_2
XFILLER_32_624 VPWR VGND sg13g2_decap_4
XFILLER_32_679 VPWR VGND sg13g2_fill_1
X_2740_ u_usb_cdc.endp\[3\] _1985_ _0984_ _0987_ _0988_ VPWR VGND sg13g2_nor4_1
X_2671_ VPWR _0940_ _0939_ VGND sg13g2_inv_1
X_4410_ net731 VGND VPWR net388 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_2
X_4341_ net686 VGND VPWR _0343_ u_usb_cdc.u_sie.data_q\[4\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4272_ net680 VGND VPWR _0274_ u_usb_cdc.addr\[6\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
X_3223_ VPWR VGND _1279_ _1293_ _1290_ net808 _1294_ _1289_ sg13g2_a221oi_1
X_3154_ _1234_ VPWR _0234_ VGND _1173_ _1229_ sg13g2_o21ai_1
XFILLER_28_908 VPWR VGND sg13g2_fill_1
X_3085_ _1197_ VPWR _0202_ VGND net719 net607 sg13g2_o21ai_1
X_2105_ VPWR _1983_ net136 VGND sg13g2_inv_1
X_2036_ net786 _1915_ VPWR VGND sg13g2_inv_4
XFILLER_36_996 VPWR VGND sg13g2_decap_8
X_3987_ _2001_ net1000 _1871_ VPWR VGND sg13g2_xor2_1
XFILLER_11_808 VPWR VGND sg13g2_fill_2
XFILLER_22_145 VPWR VGND sg13g2_fill_1
X_2938_ _1116_ VPWR _0136_ VGND net707 _1093_ sg13g2_o21ai_1
X_2869_ _1084_ net89 _1080_ VPWR VGND sg13g2_nand2_1
Xhold330 u_usb_cdc.u_sie.crc16_q\[3\] VPWR VGND net372 sg13g2_dlygate4sd3_1
Xhold352 _0390_ VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold341 _0037_ VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold385 _0109_ VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold396 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[7\] VPWR VGND
+ net438 sg13g2_dlygate4sd3_1
Xhold363 _1276_ VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold374 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[49\] VPWR
+ VGND net416 sg13g2_dlygate4sd3_1
Xfanout810 net811 net810 VPWR VGND sg13g2_buf_8
Xfanout821 net1057 net821 VPWR VGND sg13g2_buf_8
Xfanout832 net981 net832 VPWR VGND sg13g2_buf_8
XFILLER_19_919 VPWR VGND sg13g2_fill_1
XFILLER_42_900 VPWR VGND sg13g2_decap_8
XFILLER_27_985 VPWR VGND sg13g2_fill_1
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_977 VPWR VGND sg13g2_decap_8
XFILLER_41_487 VPWR VGND sg13g2_decap_8
XFILLER_13_189 VPWR VGND sg13g2_fill_1
XFILLER_5_311 VPWR VGND sg13g2_fill_1
XFILLER_6_856 VPWR VGND sg13g2_decap_8
XFILLER_5_388 VPWR VGND sg13g2_decap_8
XFILLER_1_561 VPWR VGND sg13g2_decap_8
XFILLER_3_68 VPWR VGND sg13g2_fill_1
XFILLER_49_554 VPWR VGND sg13g2_decap_8
XFILLER_49_598 VPWR VGND sg13g2_decap_4
XFILLER_18_930 VPWR VGND sg13g2_decap_8
XFILLER_17_451 VPWR VGND sg13g2_fill_1
XFILLER_33_911 VPWR VGND sg13g2_decap_4
X_3910_ VGND VPWR net735 _0952_ _0420_ net235 sg13g2_a21oi_1
XFILLER_33_944 VPWR VGND sg13g2_decap_8
X_3841_ _1739_ VPWR _1766_ VGND net393 _1762_ sg13g2_o21ai_1
X_3772_ _0589_ _0591_ _0981_ _1715_ _1716_ VPWR VGND sg13g2_nor4_1
XFILLER_32_487 VPWR VGND sg13g2_fill_1
X_2723_ net741 net520 _0043_ VPWR VGND sg13g2_nor2_1
XFILLER_8_193 VPWR VGND sg13g2_decap_8
X_2654_ _0925_ net892 net703 VPWR VGND sg13g2_nand2_1
X_2585_ _0646_ net888 _0867_ _0017_ VPWR VGND sg13g2_a21o_1
X_4324_ net688 VGND VPWR _0326_ u_usb_cdc.u_sie.crc16_q\[3\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_41_1003 VPWR VGND sg13g2_decap_8
X_4255_ net642 VGND VPWR net1025 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[2\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_2
X_3206_ _1278_ net811 VPWR VGND net808 sg13g2_nand2b_2
X_4186_ net645 VGND VPWR net268 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[22\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_28_716 VPWR VGND sg13g2_fill_2
X_3137_ _1225_ net248 net627 VPWR VGND sg13g2_nand2_1
XFILLER_27_204 VPWR VGND sg13g2_fill_2
X_3068_ _1188_ VPWR _0194_ VGND net719 net610 sg13g2_o21ai_1
XFILLER_36_760 VPWR VGND sg13g2_decap_4
X_2019_ _1898_ net753 VPWR VGND sg13g2_inv_8
XFILLER_3_815 VPWR VGND sg13g2_decap_8
Xhold160 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[2\] VPWR VGND net202 sg13g2_dlygate4sd3_1
Xhold171 u_usb_cdc.u_sie.addr_q\[2\] VPWR VGND net213 sg13g2_dlygate4sd3_1
Xhold182 _0223_ VPWR VGND net224 sg13g2_dlygate4sd3_1
Xhold193 _1804_ VPWR VGND net235 sg13g2_dlygate4sd3_1
Xfanout640 net643 net640 VPWR VGND sg13g2_buf_8
Xfanout651 net652 net651 VPWR VGND sg13g2_buf_8
Xfanout662 net664 net662 VPWR VGND sg13g2_buf_8
Xfanout673 net675 net673 VPWR VGND sg13g2_buf_2
Xfanout684 net685 net684 VPWR VGND sg13g2_buf_8
Xfanout695 net697 net695 VPWR VGND sg13g2_buf_8
XFILLER_37_96 VPWR VGND sg13g2_decap_8
XFILLER_14_443 VPWR VGND sg13g2_fill_1
XFILLER_10_682 VPWR VGND sg13g2_fill_1
X_2370_ _0670_ net776 VPWR VGND net774 sg13g2_nand2b_2
XFILLER_49_351 VPWR VGND sg13g2_fill_1
XFILLER_49_340 VPWR VGND sg13g2_fill_2
X_4040_ net678 VGND VPWR net948 u_usb_cdc.ctrl_stall clknet_leaf_48_clk sg13g2_dfrbpq_2
XFILLER_49_384 VPWR VGND sg13g2_fill_1
XFILLER_45_590 VPWR VGND sg13g2_fill_2
XFILLER_20_402 VPWR VGND sg13g2_decap_8
XFILLER_21_925 VPWR VGND sg13g2_decap_8
X_3824_ _1753_ net278 net287 _1747_ VPWR VGND sg13g2_and3_2
X_3755_ net839 VPWR _1701_ VGND _0579_ _1018_ sg13g2_o21ai_1
X_3686_ net794 VPWR _1656_ VGND net802 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[54\]
+ sg13g2_o21ai_1
XFILLER_9_491 VPWR VGND sg13g2_decap_8
X_2706_ _0964_ net807 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[2\]
+ VPWR VGND sg13g2_xnor2_1
X_2637_ _0529_ _0908_ _0909_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_829 VPWR VGND sg13g2_decap_8
X_2568_ VPWR _0012_ net1038 VGND sg13g2_inv_1
X_2499_ VPWR VGND _0795_ _0793_ _0794_ net760 _0796_ net758 sg13g2_a221oi_1
X_4307_ net679 VGND VPWR _0309_ u_usb_cdc.u_sie.addr_q\[3\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_4238_ net646 VGND VPWR net1058 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[2\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_2
XFILLER_28_524 VPWR VGND sg13g2_decap_8
X_4169_ net663 VGND VPWR net233 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[5\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_11_457 VPWR VGND sg13g2_decap_4
XFILLER_12_958 VPWR VGND sg13g2_decap_8
XFILLER_3_689 VPWR VGND sg13g2_decap_8
XFILLER_2_155 VPWR VGND sg13g2_fill_1
XFILLER_47_800 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_47_877 VPWR VGND sg13g2_decap_8
XFILLER_46_398 VPWR VGND sg13g2_fill_2
XFILLER_46_387 VPWR VGND sg13g2_decap_8
XFILLER_30_700 VPWR VGND sg13g2_fill_2
XFILLER_31_1024 VPWR VGND sg13g2_decap_4
XFILLER_7_962 VPWR VGND sg13g2_decap_8
XFILLER_11_980 VPWR VGND sg13g2_decap_8
X_3540_ _1516_ _1917_ u_usb_cdc.u_ctrl_endp.req_q\[8\] VPWR VGND sg13g2_nand2_2
XFILLER_6_461 VPWR VGND sg13g2_fill_1
X_3471_ _1468_ _1469_ _0316_ VPWR VGND sg13g2_nor2_1
X_2422_ _0718_ _0719_ _0716_ _0720_ VPWR VGND sg13g2_nand3_1
X_2353_ net779 _0649_ _0653_ VPWR VGND sg13g2_nor2_2
X_4023_ net667 VGND VPWR net954 u_usb_cdc.u_ctrl_endp.req_q\[3\] clknet_leaf_49_clk
+ sg13g2_dfrbpq_1
X_2284_ _0586_ _0053_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] VPWR VGND sg13g2_nand2b_1
XFILLER_38_822 VPWR VGND sg13g2_decap_4
XFILLER_49_192 VPWR VGND sg13g2_decap_4
XFILLER_49_170 VPWR VGND sg13g2_fill_2
XFILLER_37_321 VPWR VGND sg13g2_decap_4
XFILLER_25_505 VPWR VGND sg13g2_fill_2
XFILLER_38_877 VPWR VGND sg13g2_decap_8
XFILLER_37_387 VPWR VGND sg13g2_decap_4
X_3807_ net318 net600 _1741_ VPWR VGND sg13g2_nor2_1
X_3738_ net752 net503 _0602_ _0361_ VPWR VGND sg13g2_mux2_1
X_3669_ VPWR VGND _1639_ _1516_ _1617_ _0552_ _1640_ _0850_ sg13g2_a221oi_1
XFILLER_0_626 VPWR VGND sg13g2_decap_8
XFILLER_44_836 VPWR VGND sg13g2_decap_8
XFILLER_28_387 VPWR VGND sg13g2_fill_1
XFILLER_34_42 VPWR VGND sg13g2_decap_8
XFILLER_15_1019 VPWR VGND sg13g2_decap_8
XFILLER_11_265 VPWR VGND sg13g2_decap_4
XFILLER_8_748 VPWR VGND sg13g2_decap_8
XFILLER_4_921 VPWR VGND sg13g2_decap_8
XFILLER_4_998 VPWR VGND sg13g2_decap_8
XFILLER_43_880 VPWR VGND sg13g2_decap_8
X_2971_ VPWR _0158_ _1127_ VGND sg13g2_inv_1
Xhold737 _0255_ VPWR VGND net1055 sg13g2_dlygate4sd3_1
Xhold726 u_usb_cdc.sie_out_err VPWR VGND net1044 sg13g2_dlygate4sd3_1
Xhold715 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ VPWR VGND net1033 sg13g2_dlygate4sd3_1
Xhold704 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ VPWR VGND net1022 sg13g2_dlygate4sd3_1
X_3523_ VGND VPWR _1496_ _1498_ _1499_ net788 sg13g2_a21oi_1
Xhold748 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[1\] VPWR VGND
+ net1066 sg13g2_dlygate4sd3_1
XFILLER_6_291 VPWR VGND sg13g2_fill_1
X_3454_ _1456_ _0647_ _1455_ net878 net738 VPWR VGND sg13g2_a22oi_1
X_2405_ net784 _0661_ _0705_ VPWR VGND sg13g2_nor2_2
X_3385_ net757 _1408_ _1411_ VPWR VGND sg13g2_nor2_1
X_2336_ _0635_ net738 _0637_ VPWR VGND _0631_ sg13g2_nand3b_1
X_2267_ _0564_ _0565_ net767 _0569_ VPWR VGND _0566_ sg13g2_nand4_1
Xclkbuf_leaf_49_clk clknet_3_1__leaf_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
XFILLER_29_129 VPWR VGND sg13g2_fill_2
X_4006_ _1885_ net632 _1884_ VPWR VGND sg13g2_nand2_1
X_2198_ u_usb_cdc.u_sie.data_q\[7\] net881 _0500_ VPWR VGND sg13g2_xor2_1
XFILLER_38_1019 VPWR VGND sg13g2_decap_4
XFILLER_5_729 VPWR VGND sg13g2_decap_8
XFILLER_0_423 VPWR VGND sg13g2_decap_8
XFILLER_1_946 VPWR VGND sg13g2_decap_8
XFILLER_49_928 VPWR VGND sg13g2_decap_8
Xhold20 _0103_ VPWR VGND net62 sg13g2_dlygate4sd3_1
Xhold31 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[41\] VPWR VGND
+ net73 sg13g2_dlygate4sd3_1
XFILLER_48_449 VPWR VGND sg13g2_fill_2
Xhold64 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[53\] VPWR VGND
+ net106 sg13g2_dlygate4sd3_1
Xhold53 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[8\] VPWR VGND
+ net95 sg13g2_dlygate4sd3_1
Xhold42 _0123_ VPWR VGND net84 sg13g2_dlygate4sd3_1
Xhold97 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[38\] VPWR VGND
+ net139 sg13g2_dlygate4sd3_1
Xhold75 _0237_ VPWR VGND net117 sg13g2_dlygate4sd3_1
Xhold86 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[62\] VPWR VGND
+ net128 sg13g2_dlygate4sd3_1
XFILLER_21_1012 VPWR VGND sg13g2_decap_8
XFILLER_21_1023 VPWR VGND sg13g2_fill_2
XFILLER_29_696 VPWR VGND sg13g2_decap_4
XFILLER_40_850 VPWR VGND sg13g2_fill_1
XFILLER_4_795 VPWR VGND sg13g2_decap_8
XFILLER_3_272 VPWR VGND sg13g2_fill_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_1017 VPWR VGND sg13g2_decap_8
X_3170_ _1246_ net807 _1245_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_405 VPWR VGND sg13g2_fill_2
XFILLER_0_990 VPWR VGND sg13g2_decap_8
X_2121_ _1999_ net743 _1997_ VPWR VGND sg13g2_nand2_2
X_2052_ VPWR _1931_ u_usb_cdc.u_ctrl_endp.req_q\[6\] VGND sg13g2_inv_1
XFILLER_48_994 VPWR VGND sg13g2_decap_8
XFILLER_31_850 VPWR VGND sg13g2_fill_2
X_2954_ net450 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ _1121_ _0147_ VPWR VGND sg13g2_mux2_1
X_2885_ _1095_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ _1082_ VPWR VGND sg13g2_nand2_1
Xhold501 _0074_ VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold512 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[5\] VPWR VGND
+ net554 sg13g2_dlygate4sd3_1
X_3506_ _0335_ net572 _1951_ net575 _1941_ VPWR VGND sg13g2_a22oi_1
Xhold534 u_usb_cdc.u_sie.u_phy_rx.dp_q\[0\] VPWR VGND net852 sg13g2_dlygate4sd3_1
Xhold545 _1726_ VPWR VGND net863 sg13g2_dlygate4sd3_1
Xhold523 _1892_ VPWR VGND net565 sg13g2_dlygate4sd3_1
Xhold567 _0286_ VPWR VGND net885 sg13g2_dlygate4sd3_1
Xhold578 u_usb_cdc.addr\[4\] VPWR VGND net896 sg13g2_dlygate4sd3_1
Xhold556 net36 VPWR VGND net874 sg13g2_dlygate4sd3_1
Xhold589 _0007_ VPWR VGND net907 sg13g2_dlygate4sd3_1
X_3437_ VGND VPWR _1907_ net582 _0304_ _1447_ sg13g2_a21oi_1
X_3368_ _0724_ _1398_ _1399_ VPWR VGND sg13g2_nor2_2
X_2319_ _0588_ VPWR _0620_ VGND _0613_ _0619_ sg13g2_o21ai_1
X_3299_ _0257_ net808 _1354_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_471 VPWR VGND sg13g2_decap_8
XFILLER_39_994 VPWR VGND sg13g2_decap_8
XFILLER_25_132 VPWR VGND sg13g2_decap_8
XFILLER_26_644 VPWR VGND sg13g2_decap_8
XFILLER_25_154 VPWR VGND sg13g2_decap_8
XFILLER_26_699 VPWR VGND sg13g2_decap_8
XFILLER_41_636 VPWR VGND sg13g2_decap_8
XFILLER_40_146 VPWR VGND sg13g2_fill_2
XFILLER_5_537 VPWR VGND sg13g2_decap_4
XFILLER_31_87 VPWR VGND sg13g2_fill_2
Xoutput32 net32 uo_out[3] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uio_oe[7] VPWR VGND sg13g2_buf_1
XFILLER_0_220 VPWR VGND sg13g2_fill_2
XFILLER_1_743 VPWR VGND sg13g2_decap_8
XFILLER_49_725 VPWR VGND sg13g2_decap_8
XFILLER_0_286 VPWR VGND sg13g2_decap_8
XFILLER_17_600 VPWR VGND sg13g2_fill_2
XFILLER_36_419 VPWR VGND sg13g2_fill_2
XFILLER_45_975 VPWR VGND sg13g2_decap_8
X_2670_ _0915_ _0919_ net935 _0939_ VPWR VGND _0936_ sg13g2_nand4_1
X_4340_ net686 VGND VPWR _0342_ u_usb_cdc.u_sie.data_q\[3\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4271_ net693 VGND VPWR _0273_ u_usb_cdc.addr\[5\] clknet_leaf_43_clk sg13g2_dfrbpq_2
X_3222_ _1278_ _1291_ _1292_ _1293_ VPWR VGND sg13g2_nor3_1
X_3153_ _1234_ net193 _1230_ VPWR VGND sg13g2_nand2_1
X_2104_ VPWR _1982_ net860 VGND sg13g2_inv_1
XFILLER_27_408 VPWR VGND sg13g2_decap_8
XFILLER_48_791 VPWR VGND sg13g2_decap_8
X_3084_ _1197_ net77 net607 VPWR VGND sg13g2_nand2_1
X_2035_ _1914_ net788 VPWR VGND sg13g2_inv_2
XFILLER_36_975 VPWR VGND sg13g2_decap_8
XFILLER_22_113 VPWR VGND sg13g2_decap_4
X_3986_ VGND VPWR _1998_ _1870_ _0430_ _1869_ sg13g2_a21oi_1
X_2937_ _1116_ net106 _1110_ VPWR VGND sg13g2_nand2_1
XFILLER_11_1022 VPWR VGND sg13g2_decap_8
X_2868_ _1081_ VPWR _0099_ VGND net826 _1083_ sg13g2_o21ai_1
X_2799_ net828 net827 net824 _1040_ VPWR VGND sg13g2_nor3_2
Xhold320 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[48\] VPWR
+ VGND net362 sg13g2_dlygate4sd3_1
Xhold331 _0334_ VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold342 u_usb_cdc.u_ctrl_endp.addr_dd\[4\] VPWR VGND net384 sg13g2_dlygate4sd3_1
XFILLER_2_529 VPWR VGND sg13g2_decap_8
Xhold353 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[56\] VPWR VGND
+ net395 sg13g2_dlygate4sd3_1
Xfanout800 net804 net800 VPWR VGND sg13g2_buf_8
Xhold364 _0243_ VPWR VGND net406 sg13g2_dlygate4sd3_1
Xhold375 _0216_ VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold386 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[5\] VPWR VGND net428 sg13g2_dlygate4sd3_1
Xhold397 _0090_ VPWR VGND net439 sg13g2_dlygate4sd3_1
Xfanout811 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[1\] net811
+ VPWR VGND sg13g2_buf_8
Xfanout822 net823 net822 VPWR VGND sg13g2_buf_8
Xfanout833 net847 net833 VPWR VGND sg13g2_buf_8
XFILLER_46_739 VPWR VGND sg13g2_decap_8
XFILLER_26_43 VPWR VGND sg13g2_fill_2
XFILLER_42_956 VPWR VGND sg13g2_decap_8
XFILLER_13_135 VPWR VGND sg13g2_fill_2
XFILLER_6_835 VPWR VGND sg13g2_decap_8
XFILLER_5_367 VPWR VGND sg13g2_decap_8
XFILLER_3_47 VPWR VGND sg13g2_decap_4
XFILLER_1_540 VPWR VGND sg13g2_decap_8
XFILLER_49_533 VPWR VGND sg13g2_decap_8
XFILLER_45_783 VPWR VGND sg13g2_decap_8
XFILLER_45_750 VPWR VGND sg13g2_decap_8
XFILLER_17_463 VPWR VGND sg13g2_decap_8
XFILLER_32_411 VPWR VGND sg13g2_fill_2
X_3840_ net393 _1762_ _1765_ VPWR VGND sg13g2_and2_1
XFILLER_20_617 VPWR VGND sg13g2_decap_8
X_3771_ _1715_ _1714_ _0494_ _1706_ _0908_ VPWR VGND sg13g2_a22oi_1
XFILLER_34_1022 VPWR VGND sg13g2_decap_8
X_2722_ net519 _0454_ _0975_ VPWR VGND sg13g2_nor2_1
X_2653_ net635 _0453_ net257 _0924_ VPWR VGND sg13g2_nand3_1
X_2584_ _0639_ _0640_ _0866_ _0867_ VPWR VGND sg13g2_nor3_1
X_4323_ net688 VGND VPWR _0325_ u_usb_cdc.u_sie.crc16_q\[2\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_5_890 VPWR VGND sg13g2_decap_8
X_4254_ net642 VGND VPWR _0256_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[1\]
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3205_ net815 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[32\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[40\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[48\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[56\] net811 _1277_
+ VPWR VGND sg13g2_mux4_1
X_4185_ net646 VGND VPWR net284 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[21\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3136_ _1224_ VPWR _0226_ VGND net719 net629 sg13g2_o21ai_1
X_3067_ _1188_ net58 net610 VPWR VGND sg13g2_nand2_1
X_2018_ VPWR _1897_ net756 VGND sg13g2_inv_1
XFILLER_23_455 VPWR VGND sg13g2_decap_4
XFILLER_24_989 VPWR VGND sg13g2_decap_8
XFILLER_10_149 VPWR VGND sg13g2_decap_8
X_3969_ _1857_ _1947_ net831 _1924_ net830 VPWR VGND sg13g2_a22oi_1
Xhold150 _0093_ VPWR VGND net192 sg13g2_dlygate4sd3_1
Xhold161 _0383_ VPWR VGND net203 sg13g2_dlygate4sd3_1
Xhold172 u_usb_cdc.u_sie.addr_q\[5\] VPWR VGND net214 sg13g2_dlygate4sd3_1
Xhold194 _0420_ VPWR VGND net236 sg13g2_dlygate4sd3_1
Xhold183 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[13\] VPWR
+ VGND net225 sg13g2_dlygate4sd3_1
Xfanout630 _1135_ net630 VPWR VGND sg13g2_buf_8
Xfanout641 net642 net641 VPWR VGND sg13g2_buf_8
Xfanout663 net664 net663 VPWR VGND sg13g2_buf_8
Xfanout652 net658 net652 VPWR VGND sg13g2_buf_8
Xfanout685 net690 net685 VPWR VGND sg13g2_buf_8
Xfanout674 net675 net674 VPWR VGND sg13g2_buf_8
XFILLER_19_739 VPWR VGND sg13g2_fill_1
Xfanout696 net697 net696 VPWR VGND sg13g2_buf_8
XFILLER_37_31 VPWR VGND sg13g2_fill_2
XFILLER_37_75 VPWR VGND sg13g2_fill_1
XFILLER_14_411 VPWR VGND sg13g2_decap_8
XFILLER_15_934 VPWR VGND sg13g2_fill_2
XFILLER_26_260 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_131 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_4
XFILLER_2_893 VPWR VGND sg13g2_decap_8
XFILLER_37_536 VPWR VGND sg13g2_decap_4
X_3823_ _1751_ VPWR _0385_ VGND net278 _1752_ sg13g2_o21ai_1
XFILLER_20_414 VPWR VGND sg13g2_fill_2
X_3754_ net1009 _1700_ _1695_ _0368_ VPWR VGND sg13g2_mux2_1
X_3685_ _1912_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[62\] _1655_
+ VPWR VGND sg13g2_nor2_1
X_2705_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[3\] net806
+ _0963_ VPWR VGND sg13g2_xor2_1
X_2636_ net745 _1903_ _0908_ VPWR VGND sg13g2_nor2_1
XFILLER_0_808 VPWR VGND sg13g2_decap_8
X_2567_ VPWR VGND net739 _0854_ _0695_ net1037 _0855_ _0646_ sg13g2_a221oi_1
X_2498_ _0480_ _0730_ _0795_ VPWR VGND sg13g2_nor2_1
X_4306_ net693 VGND VPWR _0308_ u_usb_cdc.u_sie.addr_q\[2\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_4237_ net646 VGND VPWR _0240_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\]
+ clknet_leaf_4_clk sg13g2_dfrbpq_2
XFILLER_28_503 VPWR VGND sg13g2_fill_2
X_4168_ net661 VGND VPWR net158 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[4\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_4099_ net651 VGND VPWR net185 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[19\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3119_ VGND VPWR _1173_ net604 _0218_ _1215_ sg13g2_a21oi_1
XFILLER_16_709 VPWR VGND sg13g2_fill_1
XFILLER_12_937 VPWR VGND sg13g2_decap_8
XFILLER_23_274 VPWR VGND sg13g2_fill_1
XFILLER_11_436 VPWR VGND sg13g2_fill_1
XFILLER_3_668 VPWR VGND sg13g2_decap_8
XFILLER_24_1010 VPWR VGND sg13g2_decap_8
XFILLER_47_856 VPWR VGND sg13g2_decap_8
XFILLER_14_230 VPWR VGND sg13g2_fill_2
XFILLER_30_767 VPWR VGND sg13g2_fill_1
XFILLER_31_1003 VPWR VGND sg13g2_decap_8
XFILLER_7_941 VPWR VGND sg13g2_decap_8
X_3470_ _1467_ VPWR _1469_ VGND net1005 net742 sg13g2_o21ai_1
X_2421_ net617 VPWR _0719_ VGND _0694_ _0696_ sg13g2_o21ai_1
XFILLER_9_1015 VPWR VGND sg13g2_decap_8
X_2352_ net715 _0650_ net786 _0652_ VPWR VGND sg13g2_nand3_1
XFILLER_2_690 VPWR VGND sg13g2_decap_8
X_2283_ _0585_ _1993_ net705 VPWR VGND sg13g2_nand2_2
X_4022_ net666 VGND VPWR _0003_ u_usb_cdc.u_ctrl_endp.req_q\[2\] clknet_leaf_49_clk
+ sg13g2_dfrbpq_2
XFILLER_37_300 VPWR VGND sg13g2_decap_8
X_3806_ _1740_ net740 VPWR VGND _1738_ sg13g2_nand2b_2
X_3737_ net753 net370 net589 _0360_ VPWR VGND sg13g2_mux2_1
X_3668_ _1639_ _1519_ net773 VPWR VGND sg13g2_nand2b_1
XFILLER_47_1010 VPWR VGND sg13g2_decap_8
X_3599_ _0542_ _0670_ _1573_ VPWR VGND sg13g2_nor2_1
X_2619_ VGND VPWR net838 net593 _0898_ _0897_ sg13g2_a21oi_1
XFILLER_0_605 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_fill_2
XFILLER_28_322 VPWR VGND sg13g2_fill_1
XFILLER_44_815 VPWR VGND sg13g2_decap_8
XFILLER_28_344 VPWR VGND sg13g2_decap_8
XFILLER_28_366 VPWR VGND sg13g2_fill_1
XFILLER_24_561 VPWR VGND sg13g2_decap_8
XFILLER_8_738 VPWR VGND sg13g2_decap_4
XFILLER_4_900 VPWR VGND sg13g2_decap_8
XFILLER_4_977 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_15_8 VPWR VGND sg13g2_fill_2
XFILLER_35_859 VPWR VGND sg13g2_fill_1
X_2970_ net638 VPWR _1127_ VGND net941 _1056_ sg13g2_o21ai_1
XFILLER_34_369 VPWR VGND sg13g2_decap_8
XFILLER_30_564 VPWR VGND sg13g2_decap_8
XFILLER_30_575 VPWR VGND sg13g2_fill_2
XFILLER_7_782 VPWR VGND sg13g2_decap_8
Xhold716 u_usb_cdc.sie_in_data_ack VPWR VGND net1034 sg13g2_dlygate4sd3_1
Xhold705 u_usb_cdc.u_sie.data_q\[2\] VPWR VGND net1023 sg13g2_dlygate4sd3_1
X_3522_ VGND VPWR net792 _1497_ _1498_ _1913_ sg13g2_a21oi_1
Xhold727 u_usb_cdc.u_sie.phy_state_q\[7\] VPWR VGND net1045 sg13g2_dlygate4sd3_1
Xhold749 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[0\] VPWR VGND
+ net1067 sg13g2_dlygate4sd3_1
X_3453_ VGND VPWR _1932_ _1383_ _1455_ _0614_ sg13g2_a21oi_1
Xhold738 u_usb_cdc.bulk_out_nak[0] VPWR VGND net1056 sg13g2_dlygate4sd3_1
X_2404_ _1901_ _0478_ _1899_ _0704_ VPWR VGND _0702_ sg13g2_nand4_1
X_3384_ net856 net567 _1410_ VPWR VGND sg13g2_nor2_1
X_2335_ _0636_ _0635_ _0631_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_631 VPWR VGND sg13g2_fill_1
X_2266_ _0567_ VPWR _0568_ VGND _1914_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\]
+ sg13g2_o21ai_1
XFILLER_26_804 VPWR VGND sg13g2_fill_2
X_2197_ net832 VPWR _0499_ VGND _0469_ _0498_ sg13g2_o21ai_1
X_4005_ net594 _1883_ _1884_ VPWR VGND sg13g2_nor2_1
XFILLER_26_848 VPWR VGND sg13g2_fill_2
XFILLER_38_686 VPWR VGND sg13g2_fill_2
XFILLER_25_336 VPWR VGND sg13g2_decap_4
XFILLER_25_358 VPWR VGND sg13g2_fill_2
XFILLER_37_196 VPWR VGND sg13g2_decap_8
XFILLER_41_818 VPWR VGND sg13g2_decap_8
XFILLER_33_380 VPWR VGND sg13g2_decap_8
XFILLER_34_892 VPWR VGND sg13g2_fill_2
XFILLER_21_575 VPWR VGND sg13g2_decap_4
XFILLER_5_708 VPWR VGND sg13g2_decap_8
XFILLER_0_402 VPWR VGND sg13g2_decap_8
XFILLER_1_925 VPWR VGND sg13g2_decap_8
XFILLER_49_907 VPWR VGND sg13g2_decap_8
Xhold21 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[3\] VPWR VGND
+ net63 sg13g2_dlygate4sd3_1
XFILLER_0_479 VPWR VGND sg13g2_decap_8
Xhold10 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[2\] VPWR VGND net52 sg13g2_dlygate4sd3_1
Xhold32 _0124_ VPWR VGND net74 sg13g2_dlygate4sd3_1
Xhold65 _0136_ VPWR VGND net107 sg13g2_dlygate4sd3_1
Xhold54 _0091_ VPWR VGND net96 sg13g2_dlygate4sd3_1
XFILLER_29_54 VPWR VGND sg13g2_decap_8
XFILLER_29_631 VPWR VGND sg13g2_decap_8
Xhold43 u_usb_cdc.u_sie.in_zlp_q\[1\] VPWR VGND net85 sg13g2_dlygate4sd3_1
Xhold98 _0205_ VPWR VGND net140 sg13g2_dlygate4sd3_1
Xhold76 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[64\] VPWR VGND
+ net118 sg13g2_dlygate4sd3_1
Xhold87 _0229_ VPWR VGND net129 sg13g2_dlygate4sd3_1
XFILLER_43_111 VPWR VGND sg13g2_fill_1
XFILLER_24_380 VPWR VGND sg13g2_decap_4
XFILLER_8_524 VPWR VGND sg13g2_fill_2
XFILLER_4_774 VPWR VGND sg13g2_decap_8
XFILLER_3_251 VPWR VGND sg13g2_fill_2
X_2120_ net713 _1996_ _1998_ VPWR VGND sg13g2_nor2_1
XFILLER_48_973 VPWR VGND sg13g2_decap_8
X_2051_ VPWR _1930_ net868 VGND sg13g2_inv_1
XFILLER_19_130 VPWR VGND sg13g2_decap_4
XFILLER_47_494 VPWR VGND sg13g2_decap_8
XFILLER_34_122 VPWR VGND sg13g2_fill_1
X_2953_ _1121_ net736 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ _1040_ VPWR VGND sg13g2_and3_2
XFILLER_22_339 VPWR VGND sg13g2_fill_2
X_2884_ _1094_ net147 _1080_ VPWR VGND sg13g2_nand2_1
XFILLER_30_372 VPWR VGND sg13g2_decap_4
Xhold502 net33 VPWR VGND net544 sg13g2_dlygate4sd3_1
Xhold513 _0088_ VPWR VGND net555 sg13g2_dlygate4sd3_1
X_3505_ _0334_ net572 _1948_ net577 _1942_ VPWR VGND sg13g2_a22oi_1
Xhold524 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] VPWR VGND net566 sg13g2_dlygate4sd3_1
Xhold535 _0409_ VPWR VGND net853 sg13g2_dlygate4sd3_1
Xhold568 u_usb_cdc.addr\[6\] VPWR VGND net886 sg13g2_dlygate4sd3_1
Xhold557 _0250_ VPWR VGND net875 sg13g2_dlygate4sd3_1
Xhold579 net34 VPWR VGND net897 sg13g2_dlygate4sd3_1
Xhold546 u_usb_cdc.u_ctrl_endp.max_length_q\[0\] VPWR VGND net864 sg13g2_dlygate4sd3_1
X_3436_ net766 net582 _1447_ VPWR VGND sg13g2_nor2_1
X_3367_ VGND VPWR _0653_ _0705_ _1398_ net620 sg13g2_a21oi_1
X_2318_ _0563_ _0570_ _0615_ _0618_ _0619_ VPWR VGND sg13g2_nor4_1
X_3298_ net809 net807 net812 _1356_ VPWR VGND _1274_ sg13g2_nand4_1
XFILLER_39_973 VPWR VGND sg13g2_decap_8
X_2249_ net780 net777 _0549_ _0551_ VPWR VGND sg13g2_nor3_2
XFILLER_25_111 VPWR VGND sg13g2_fill_1
XFILLER_13_328 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_fill_2
Xoutput33 net33 uo_out[4] VPWR VGND sg13g2_buf_1
Xoutput22 net22 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_722 VPWR VGND sg13g2_decap_8
XFILLER_49_704 VPWR VGND sg13g2_decap_8
XFILLER_1_799 VPWR VGND sg13g2_decap_8
XFILLER_0_298 VPWR VGND sg13g2_decap_8
XFILLER_45_954 VPWR VGND sg13g2_decap_8
XFILLER_17_678 VPWR VGND sg13g2_fill_1
XFILLER_32_659 VPWR VGND sg13g2_fill_2
XFILLER_9_866 VPWR VGND sg13g2_decap_8
X_4270_ net693 VGND VPWR _0272_ u_usb_cdc.addr\[4\] clknet_leaf_43_clk sg13g2_dfrbpq_2
XFILLER_28_1019 VPWR VGND sg13g2_decap_8
X_3221_ net815 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[17\]
+ _1292_ VPWR VGND sg13g2_nor2_1
X_3152_ _1233_ VPWR _0233_ VGND _1172_ _1229_ sg13g2_o21ai_1
X_2103_ VPWR _1981_ net287 VGND sg13g2_inv_1
XFILLER_48_770 VPWR VGND sg13g2_decap_8
X_3083_ _1196_ VPWR _0201_ VGND net718 net606 sg13g2_o21ai_1
X_2034_ net989 _1913_ VPWR VGND sg13g2_inv_4
XFILLER_36_954 VPWR VGND sg13g2_decap_8
XFILLER_23_637 VPWR VGND sg13g2_decap_4
XFILLER_35_486 VPWR VGND sg13g2_fill_2
XFILLER_22_136 VPWR VGND sg13g2_decap_8
X_3985_ _2001_ VPWR _1870_ VGND _1993_ _1034_ sg13g2_o21ai_1
XFILLER_22_169 VPWR VGND sg13g2_decap_4
X_2936_ _1115_ VPWR _0135_ VGND net707 _1091_ sg13g2_o21ai_1
X_2867_ _1083_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ _1082_ VPWR VGND sg13g2_nand2_1
XFILLER_11_1001 VPWR VGND sg13g2_decap_8
X_2798_ net827 net825 _1039_ VPWR VGND sg13g2_nor2_1
Xhold310 _0456_ VPWR VGND net352 sg13g2_dlygate4sd3_1
Xhold343 _0279_ VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold321 _0215_ VPWR VGND net363 sg13g2_dlygate4sd3_1
Xhold332 net16 VPWR VGND net374 sg13g2_dlygate4sd3_1
Xhold365 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[3\] VPWR VGND
+ net407 sg13g2_dlygate4sd3_1
Xhold387 _1725_ VPWR VGND net429 sg13g2_dlygate4sd3_1
Xhold354 _0139_ VPWR VGND net396 sg13g2_dlygate4sd3_1
Xhold376 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[24\] VPWR VGND
+ net418 sg13g2_dlygate4sd3_1
Xfanout801 net802 net801 VPWR VGND sg13g2_buf_8
Xhold398 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[19\] VPWR
+ VGND net440 sg13g2_dlygate4sd3_1
Xfanout812 net814 net812 VPWR VGND sg13g2_buf_8
Xfanout823 net1059 net823 VPWR VGND sg13g2_buf_8
X_3419_ _0298_ _1433_ _1435_ VPWR VGND sg13g2_nand2_1
Xfanout834 net835 net834 VPWR VGND sg13g2_buf_8
X_4399_ net725 VGND VPWR net53 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[2\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_46_718 VPWR VGND sg13g2_decap_8
XFILLER_26_464 VPWR VGND sg13g2_fill_2
XFILLER_27_976 VPWR VGND sg13g2_decap_8
XFILLER_42_935 VPWR VGND sg13g2_decap_8
XFILLER_26_475 VPWR VGND sg13g2_fill_2
XFILLER_42_21 VPWR VGND sg13g2_fill_2
XFILLER_22_692 VPWR VGND sg13g2_decap_8
XFILLER_6_814 VPWR VGND sg13g2_decap_8
XFILLER_10_876 VPWR VGND sg13g2_fill_1
XFILLER_3_15 VPWR VGND sg13g2_decap_4
XFILLER_49_512 VPWR VGND sg13g2_decap_8
XFILLER_1_596 VPWR VGND sg13g2_decap_8
XFILLER_18_965 VPWR VGND sg13g2_fill_2
XFILLER_44_283 VPWR VGND sg13g2_decap_4
XFILLER_32_434 VPWR VGND sg13g2_decap_8
XFILLER_32_456 VPWR VGND sg13g2_decap_8
XFILLER_33_979 VPWR VGND sg13g2_decap_8
XFILLER_13_670 VPWR VGND sg13g2_fill_1
X_3770_ _0466_ _1713_ _1714_ VPWR VGND sg13g2_nor2_1
XFILLER_34_1001 VPWR VGND sg13g2_decap_8
X_2721_ net741 net264 _0044_ VPWR VGND sg13g2_nor2_1
X_2652_ net635 _0922_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] _0923_ VPWR VGND sg13g2_nand3_1
X_2583_ VGND VPWR u_usb_cdc.sie_in_data_ack _0865_ _0866_ net888 sg13g2_a21oi_1
X_4322_ net695 VGND VPWR _0324_ u_usb_cdc.u_sie.crc16_q\[1\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4253_ net643 VGND VPWR net1055 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[0\]
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3204_ net404 _1274_ _1276_ VPWR VGND sg13g2_nor2_1
X_4184_ net647 VGND VPWR net300 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[20\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_28_707 VPWR VGND sg13g2_fill_2
X_3135_ _1224_ net164 net629 VPWR VGND sg13g2_nand2_1
XFILLER_27_206 VPWR VGND sg13g2_fill_1
X_3066_ _1187_ VPWR _0193_ VGND net718 net608 sg13g2_o21ai_1
XFILLER_42_209 VPWR VGND sg13g2_decap_8
X_2017_ VPWR _1896_ net755 VGND sg13g2_inv_1
XFILLER_24_924 VPWR VGND sg13g2_decap_4
XFILLER_35_272 VPWR VGND sg13g2_fill_2
XFILLER_35_283 VPWR VGND sg13g2_decap_4
XFILLER_24_968 VPWR VGND sg13g2_decap_8
X_3968_ _1851_ VPWR _0426_ VGND _1855_ _1856_ sg13g2_o21ai_1
X_2919_ _1106_ VPWR _0127_ VGND _1072_ net615 sg13g2_o21ai_1
X_3899_ _1013_ VPWR _0411_ VGND _1909_ net744 sg13g2_o21ai_1
Xhold140 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[30\] VPWR
+ VGND net182 sg13g2_dlygate4sd3_1
Xhold151 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[67\] VPWR
+ VGND net193 sg13g2_dlygate4sd3_1
Xhold162 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[29\] VPWR
+ VGND net204 sg13g2_dlygate4sd3_1
Xhold173 _0311_ VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold195 u_usb_cdc.u_sie.addr_q\[4\] VPWR VGND net237 sg13g2_dlygate4sd3_1
Xhold184 _0180_ VPWR VGND net226 sg13g2_dlygate4sd3_1
Xfanout642 net643 net642 VPWR VGND sg13g2_buf_8
Xfanout620 _0658_ net620 VPWR VGND sg13g2_buf_8
Xfanout631 net632 net631 VPWR VGND sg13g2_buf_8
Xfanout664 net667 net664 VPWR VGND sg13g2_buf_8
Xfanout653 net657 net653 VPWR VGND sg13g2_buf_8
Xfanout675 net701 net675 VPWR VGND sg13g2_buf_8
Xfanout686 net689 net686 VPWR VGND sg13g2_buf_8
Xfanout697 net700 net697 VPWR VGND sg13g2_buf_8
X_4449__42 VPWR VGND net42 sg13g2_tiehi
XFILLER_15_902 VPWR VGND sg13g2_decap_4
XFILLER_26_250 VPWR VGND sg13g2_fill_1
XFILLER_18_1007 VPWR VGND sg13g2_decap_8
XFILLER_42_798 VPWR VGND sg13g2_fill_2
XFILLER_30_949 VPWR VGND sg13g2_decap_8
XFILLER_10_651 VPWR VGND sg13g2_decap_4
XFILLER_6_622 VPWR VGND sg13g2_decap_8
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_49_320 VPWR VGND sg13g2_decap_4
XFILLER_1_393 VPWR VGND sg13g2_decap_8
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_17_283 VPWR VGND sg13g2_fill_1
XFILLER_33_765 VPWR VGND sg13g2_decap_4
X_3822_ _1752_ net600 _1747_ VPWR VGND sg13g2_nand2_1
X_3753_ _1699_ VPWR _1700_ VGND _0578_ _1692_ sg13g2_o21ai_1
X_3684_ net794 _1652_ _1653_ _1654_ VPWR VGND sg13g2_nor3_1
X_2704_ _0962_ net814 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[0\]
+ VPWR VGND sg13g2_xnor2_1
X_2635_ VPWR _0018_ _0907_ VGND sg13g2_inv_1
X_4305_ net679 VGND VPWR _0307_ u_usb_cdc.u_sie.addr_q\[1\] clknet_leaf_44_clk sg13g2_dfrbpq_1
X_2566_ net750 _0624_ _0646_ _0854_ VPWR VGND sg13g2_nor3_1
X_2497_ _1927_ u_usb_cdc.u_ctrl_endp.in_dir_q u_usb_cdc.u_ctrl_endp.rec_q\[0\] _0794_
+ VPWR VGND u_usb_cdc.configured_o sg13g2_nand4_1
X_4236_ net653 VGND VPWR _0239_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[0\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_2
X_4167_ net644 VGND VPWR _0170_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[3\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3118_ net325 net604 _1215_ VPWR VGND sg13g2_nor2_1
X_4098_ net651 VGND VPWR net179 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[18\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3049_ VGND VPWR net612 _1176_ _0187_ _1175_ sg13g2_a21oi_1
XFILLER_12_916 VPWR VGND sg13g2_decap_8
XFILLER_23_12 VPWR VGND sg13g2_fill_1
XFILLER_23_253 VPWR VGND sg13g2_decap_8
XFILLER_3_647 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_47_835 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_42_551 VPWR VGND sg13g2_decap_8
XFILLER_30_735 VPWR VGND sg13g2_fill_1
XFILLER_7_920 VPWR VGND sg13g2_decap_8
XFILLER_6_430 VPWR VGND sg13g2_decap_8
XFILLER_7_997 VPWR VGND sg13g2_decap_8
X_2420_ VPWR VGND net617 _0717_ _0698_ _0654_ _0718_ net574 sg13g2_a221oi_1
X_2351_ _0651_ net786 net715 VPWR VGND sg13g2_nand2_1
XFILLER_36_4 VPWR VGND sg13g2_fill_2
X_2282_ u_usb_cdc.u_sie.phy_state_q\[11\] net259 _0581_ _0583_ _0584_ VPWR VGND sg13g2_nor4_1
X_4021_ net677 VGND VPWR net869 u_usb_cdc.u_ctrl_endp.req_q\[1\] clknet_leaf_50_clk
+ sg13g2_dfrbpq_2
XFILLER_38_813 VPWR VGND sg13g2_fill_1
XFILLER_49_172 VPWR VGND sg13g2_fill_1
XFILLER_18_592 VPWR VGND sg13g2_fill_2
X_3805_ net710 _1738_ _1739_ VPWR VGND sg13g2_nor2_2
XFILLER_20_256 VPWR VGND sg13g2_fill_2
X_3736_ net754 net858 net589 _0359_ VPWR VGND sg13g2_mux2_1
X_3667_ _1637_ VPWR _1638_ VGND _0550_ _1524_ sg13g2_o21ai_1
X_3598_ _1570_ net774 _1572_ VPWR VGND sg13g2_nor2b_1
X_2618_ _0577_ _0617_ _0896_ _0897_ VPWR VGND sg13g2_nor3_1
X_2549_ _0000_ _0838_ _0839_ VPWR VGND sg13g2_nand2_1
X_4219_ net646 VGND VPWR net273 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[55\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_301 VPWR VGND sg13g2_fill_1
XFILLER_18_78 VPWR VGND sg13g2_fill_2
XFILLER_43_359 VPWR VGND sg13g2_decap_8
XFILLER_11_212 VPWR VGND sg13g2_decap_4
XFILLER_8_717 VPWR VGND sg13g2_decap_8
XFILLER_7_227 VPWR VGND sg13g2_decap_8
XFILLER_4_956 VPWR VGND sg13g2_decap_8
XFILLER_3_466 VPWR VGND sg13g2_decap_4
XFILLER_19_356 VPWR VGND sg13g2_fill_2
XFILLER_7_761 VPWR VGND sg13g2_decap_8
X_3521_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[48\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[56\]
+ net797 _1497_ VPWR VGND sg13g2_mux2_1
Xhold706 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[2\] VPWR
+ VGND net1024 sg13g2_dlygate4sd3_1
Xhold717 _0411_ VPWR VGND net1035 sg13g2_dlygate4sd3_1
Xhold728 u_usb_cdc.sie_in_req VPWR VGND net1046 sg13g2_dlygate4sd3_1
X_3452_ _1454_ VPWR _0312_ VGND _1901_ net580 sg13g2_o21ai_1
Xhold739 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[2\] VPWR
+ VGND net1057 sg13g2_dlygate4sd3_1
X_2403_ _0703_ _0478_ _0702_ VPWR VGND sg13g2_nand2_1
X_3383_ VGND VPWR net567 _1409_ _0288_ _1407_ sg13g2_a21oi_1
X_2334_ _0635_ _0610_ _0634_ VPWR VGND sg13g2_nand2_1
XFILLER_27_0 VPWR VGND sg13g2_decap_4
X_2265_ _0567_ _1914_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\]
+ _1912_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\] VPWR VGND
+ sg13g2_a22oi_1
X_2196_ _0498_ _0494_ _0496_ VPWR VGND sg13g2_nand2_1
X_4004_ net624 VPWR _1883_ VGND _1910_ _0612_ sg13g2_o21ai_1
XFILLER_37_153 VPWR VGND sg13g2_fill_1
XFILLER_38_676 VPWR VGND sg13g2_decap_4
XFILLER_25_348 VPWR VGND sg13g2_fill_2
XFILLER_37_186 VPWR VGND sg13g2_fill_1
X_3719_ _1685_ VPWR _0348_ VGND _1895_ net598 sg13g2_o21ai_1
XFILLER_1_904 VPWR VGND sg13g2_decap_8
Xhold22 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[44\] VPWR VGND
+ net64 sg13g2_dlygate4sd3_1
XFILLER_0_458 VPWR VGND sg13g2_decap_8
Xhold11 _0401_ VPWR VGND net53 sg13g2_dlygate4sd3_1
Xhold55 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[1\] VPWR VGND
+ net97 sg13g2_dlygate4sd3_1
Xhold44 _0436_ VPWR VGND net86 sg13g2_dlygate4sd3_1
Xhold33 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[9\] VPWR VGND
+ net75 sg13g2_dlygate4sd3_1
Xhold88 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[44\] VPWR VGND
+ net130 sg13g2_dlygate4sd3_1
Xhold77 _0231_ VPWR VGND net119 sg13g2_dlygate4sd3_1
Xhold99 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[39\] VPWR VGND
+ net141 sg13g2_dlygate4sd3_1
Xhold66 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[45\] VPWR VGND
+ net108 sg13g2_dlygate4sd3_1
XFILLER_29_665 VPWR VGND sg13g2_fill_2
XFILLER_17_827 VPWR VGND sg13g2_fill_2
XFILLER_17_838 VPWR VGND sg13g2_decap_8
XFILLER_28_175 VPWR VGND sg13g2_fill_2
XFILLER_29_687 VPWR VGND sg13g2_decap_4
XFILLER_45_32 VPWR VGND sg13g2_fill_2
XFILLER_16_326 VPWR VGND sg13g2_decap_4
XFILLER_16_348 VPWR VGND sg13g2_fill_2
XFILLER_16_359 VPWR VGND sg13g2_fill_2
XFILLER_12_510 VPWR VGND sg13g2_fill_2
XFILLER_31_318 VPWR VGND sg13g2_fill_1
XFILLER_24_392 VPWR VGND sg13g2_decap_4
XFILLER_6_26 VPWR VGND sg13g2_fill_1
XFILLER_4_753 VPWR VGND sg13g2_decap_8
XFILLER_3_263 VPWR VGND sg13g2_fill_1
XFILLER_48_952 VPWR VGND sg13g2_decap_8
X_2050_ VPWR _1929_ net741 VGND sg13g2_inv_1
XFILLER_35_624 VPWR VGND sg13g2_decap_8
XFILLER_37_1010 VPWR VGND sg13g2_decap_8
XFILLER_16_882 VPWR VGND sg13g2_fill_2
X_2952_ _1120_ VPWR _0146_ VGND _1974_ net603 sg13g2_o21ai_1
X_2883_ _1092_ VPWR _0104_ VGND net826 _1093_ sg13g2_o21ai_1
XFILLER_31_874 VPWR VGND sg13g2_fill_2
X_3504_ _0333_ net573 _1949_ net575 _1943_ VPWR VGND sg13g2_a22oi_1
Xhold503 _0247_ VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold536 u_usb_cdc.u_ctrl_endp.max_length_q\[5\] VPWR VGND net854 sg13g2_dlygate4sd3_1
Xhold525 net21 VPWR VGND net843 sg13g2_dlygate4sd3_1
Xhold514 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold547 u_usb_cdc.addr\[5\] VPWR VGND net865 sg13g2_dlygate4sd3_1
Xhold569 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[12\] VPWR VGND net887 sg13g2_dlygate4sd3_1
Xhold558 net35 VPWR VGND net876 sg13g2_dlygate4sd3_1
X_3435_ VGND VPWR _1906_ net582 _0303_ _1446_ sg13g2_a21oi_1
XFILLER_44_1025 VPWR VGND sg13g2_decap_4
X_3366_ VGND VPWR _0283_ _1397_ net345 sg13g2_or2_1
X_3297_ _1354_ _1355_ _0256_ VPWR VGND sg13g2_and2_1
X_2317_ _0618_ net839 _0578_ VPWR VGND sg13g2_nand2_1
X_2248_ net781 _0549_ _0550_ VPWR VGND sg13g2_nor2_2
XFILLER_39_952 VPWR VGND sg13g2_decap_8
X_2179_ net758 net761 _0481_ VPWR VGND sg13g2_xor2_1
XFILLER_26_657 VPWR VGND sg13g2_fill_2
XFILLER_15_46 VPWR VGND sg13g2_fill_2
XFILLER_15_79 VPWR VGND sg13g2_decap_8
XFILLER_40_148 VPWR VGND sg13g2_fill_1
XFILLER_21_362 VPWR VGND sg13g2_decap_8
Xoutput34 net34 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_701 VPWR VGND sg13g2_decap_8
Xoutput23 net23 uio_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_778 VPWR VGND sg13g2_decap_8
XFILLER_45_933 VPWR VGND sg13g2_decap_8
XFILLER_31_126 VPWR VGND sg13g2_decap_4
X_3220_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[25\] net815
+ _1291_ VPWR VGND sg13g2_nor2b_1
X_3151_ _1233_ net120 _1230_ VPWR VGND sg13g2_nand2_1
X_2102_ VPWR _1980_ net244 VGND sg13g2_inv_1
X_3082_ _1196_ net174 net606 VPWR VGND sg13g2_nand2_1
X_2033_ _1912_ net803 VPWR VGND sg13g2_inv_2
XFILLER_36_933 VPWR VGND sg13g2_decap_8
XFILLER_22_104 VPWR VGND sg13g2_fill_1
X_3984_ VGND VPWR net210 net623 _1869_ net312 sg13g2_a21oi_1
X_2935_ _1115_ net126 _1110_ VPWR VGND sg13g2_nand2_1
X_2866_ _1082_ net736 _1063_ _1079_ VPWR VGND sg13g2_and3_2
XFILLER_30_181 VPWR VGND sg13g2_decap_8
Xhold300 u_usb_cdc.u_sie.u_phy_rx.state_q\[1\] VPWR VGND net342 sg13g2_dlygate4sd3_1
Xhold311 _0064_ VPWR VGND net353 sg13g2_dlygate4sd3_1
X_2797_ _1038_ net941 net10 VPWR VGND sg13g2_nand2_1
Xhold322 u_usb_cdc.u_ctrl_endp.addr_dd\[6\] VPWR VGND net364 sg13g2_dlygate4sd3_1
XFILLER_2_509 VPWR VGND sg13g2_fill_2
Xhold344 u_usb_cdc.u_sie.u_phy_rx.dn_q\[0\] VPWR VGND net386 sg13g2_dlygate4sd3_1
Xhold333 _0357_ VPWR VGND net375 sg13g2_dlygate4sd3_1
Xhold366 _0086_ VPWR VGND net408 sg13g2_dlygate4sd3_1
Xhold377 _0107_ VPWR VGND net419 sg13g2_dlygate4sd3_1
Xhold355 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[4\] VPWR VGND
+ net397 sg13g2_dlygate4sd3_1
Xfanout802 net803 net802 VPWR VGND sg13g2_buf_8
Xfanout824 net826 net824 VPWR VGND sg13g2_buf_8
Xhold399 _0186_ VPWR VGND net441 sg13g2_dlygate4sd3_1
Xfanout813 net814 net813 VPWR VGND sg13g2_buf_1
X_4398_ net725 VGND VPWR net296 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_3418_ _1434_ _0665_ _1435_ VPWR VGND _1426_ sg13g2_nand3b_1
Xhold388 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[65\] VPWR VGND
+ net430 sg13g2_dlygate4sd3_1
X_3349_ net269 net570 _1389_ VPWR VGND sg13g2_nor2_1
Xfanout835 net1045 net835 VPWR VGND sg13g2_buf_8
XFILLER_45_229 VPWR VGND sg13g2_fill_2
XFILLER_26_421 VPWR VGND sg13g2_fill_1
XFILLER_42_914 VPWR VGND sg13g2_decap_8
XFILLER_26_432 VPWR VGND sg13g2_fill_2
XFILLER_27_999 VPWR VGND sg13g2_decap_8
XFILLER_41_435 VPWR VGND sg13g2_fill_1
XFILLER_13_137 VPWR VGND sg13g2_fill_1
XFILLER_5_303 VPWR VGND sg13g2_fill_2
XFILLER_27_1020 VPWR VGND sg13g2_decap_8
XFILLER_1_575 VPWR VGND sg13g2_decap_8
XFILLER_49_568 VPWR VGND sg13g2_fill_2
XFILLER_18_944 VPWR VGND sg13g2_fill_2
XFILLER_29_292 VPWR VGND sg13g2_fill_2
XFILLER_32_413 VPWR VGND sg13g2_fill_1
XFILLER_33_958 VPWR VGND sg13g2_decap_8
X_2720_ VGND VPWR u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[1\] net635 _0974_ net263 sg13g2_a21oi_1
XFILLER_8_163 VPWR VGND sg13g2_fill_1
X_2651_ _0919_ _0921_ _0916_ _0922_ VPWR VGND sg13g2_nand3_1
X_2582_ _1920_ _0554_ _0865_ VPWR VGND sg13g2_nor2_1
X_4321_ net695 VGND VPWR _0323_ u_usb_cdc.u_sie.crc16_q\[0\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4252_ net641 VGND VPWR net534 u_usb_cdc.out_valid_o[0] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3203_ _1275_ _0967_ _0966_ VPWR VGND sg13g2_nand2b_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
XFILLER_41_1017 VPWR VGND sg13g2_decap_8
X_4183_ net639 VGND VPWR net441 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[19\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3134_ _1223_ VPWR _0225_ VGND net718 net627 sg13g2_o21ai_1
X_3065_ _1187_ net66 net608 VPWR VGND sg13g2_nand2_1
X_2016_ net757 _1895_ VPWR VGND sg13g2_inv_4
XFILLER_35_240 VPWR VGND sg13g2_fill_2
XFILLER_35_251 VPWR VGND sg13g2_decap_8
X_3967_ _1824_ VPWR _1856_ VGND u_usb_cdc.u_sie.u_phy_tx.data_q\[6\] _1819_ sg13g2_o21ai_1
X_2918_ _1106_ net130 _1101_ VPWR VGND sg13g2_nand2_1
X_3898_ VGND VPWR _1935_ net704 _0410_ net387 sg13g2_a21oi_1
Xclkbuf_leaf_30_clk clknet_3_7__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_2849_ _1070_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net636 VPWR VGND sg13g2_nand2_1
XFILLER_3_829 VPWR VGND sg13g2_decap_8
Xhold141 _0197_ VPWR VGND net183 sg13g2_dlygate4sd3_1
Xhold152 _0234_ VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold130 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[6\] VPWR VGND net172 sg13g2_dlygate4sd3_1
Xhold174 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[9\] VPWR VGND
+ net216 sg13g2_dlygate4sd3_1
Xhold185 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[24\] VPWR
+ VGND net227 sg13g2_dlygate4sd3_1
Xhold163 _0196_ VPWR VGND net205 sg13g2_dlygate4sd3_1
Xfanout621 net622 net621 VPWR VGND sg13g2_buf_8
Xhold196 _0310_ VPWR VGND net238 sg13g2_dlygate4sd3_1
Xfanout610 _1184_ net610 VPWR VGND sg13g2_buf_8
Xfanout632 net633 net632 VPWR VGND sg13g2_buf_1
Xfanout665 net666 net665 VPWR VGND sg13g2_buf_8
Xfanout676 net677 net676 VPWR VGND sg13g2_buf_8
Xfanout643 net658 net643 VPWR VGND sg13g2_buf_8
Xfanout654 net657 net654 VPWR VGND sg13g2_buf_8
Xfanout687 net688 net687 VPWR VGND sg13g2_buf_8
Xfanout698 net700 net698 VPWR VGND sg13g2_buf_8
XFILLER_41_254 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_21_clk clknet_3_6__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_6_612 VPWR VGND sg13g2_fill_1
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_1_372 VPWR VGND sg13g2_decap_8
XFILLER_37_527 VPWR VGND sg13g2_fill_1
X_3821_ _1751_ net278 _1748_ VPWR VGND sg13g2_nand2_1
X_3752_ _0889_ _1692_ net763 _1699_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_12_clk clknet_3_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_3683_ net802 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[38\] _1653_
+ VPWR VGND sg13g2_nor2_1
X_2703_ _0961_ net810 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[1\]
+ VPWR VGND sg13g2_xnor2_1
X_2634_ _0907_ net592 net939 net596 net259 VPWR VGND sg13g2_a22oi_1
X_2565_ _0846_ VPWR _0011_ VGND _0849_ _0853_ sg13g2_o21ai_1
X_4304_ net691 VGND VPWR net965 u_usb_cdc.endp\[3\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_2496_ _0709_ _0792_ _0793_ VPWR VGND sg13g2_nor2_1
X_4235_ net643 VGND VPWR net144 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[71\]
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
X_4166_ net659 VGND VPWR _0169_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[2\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3117_ VGND VPWR _1172_ net604 _0217_ _1214_ sg13g2_a21oi_1
X_4097_ net649 VGND VPWR net90 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[17\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3048_ _1176_ net754 net630 VPWR VGND sg13g2_nand2_2
XFILLER_36_571 VPWR VGND sg13g2_fill_2
XFILLER_23_243 VPWR VGND sg13g2_fill_1
XFILLER_24_766 VPWR VGND sg13g2_fill_2
XFILLER_24_777 VPWR VGND sg13g2_fill_1
XFILLER_3_626 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_47_814 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_14_221 VPWR VGND sg13g2_decap_4
XFILLER_42_585 VPWR VGND sg13g2_decap_4
XFILLER_14_298 VPWR VGND sg13g2_fill_1
XFILLER_11_994 VPWR VGND sg13g2_decap_8
XFILLER_7_976 VPWR VGND sg13g2_decap_8
X_2350_ net777 net782 _0650_ VPWR VGND sg13g2_nor2b_2
X_2281_ VGND VPWR net208 _0582_ _0583_ net746 sg13g2_a21oi_1
X_4020_ net666 VGND VPWR net861 _0048_ clknet_leaf_50_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_29_4 VPWR VGND sg13g2_fill_2
XFILLER_38_858 VPWR VGND sg13g2_decap_4
XFILLER_18_560 VPWR VGND sg13g2_decap_8
XFILLER_21_703 VPWR VGND sg13g2_decap_4
XFILLER_33_552 VPWR VGND sg13g2_decap_4
X_3804_ net342 u_usb_cdc.u_sie.u_phy_rx.state_q\[2\] _1737_ _1738_ VPWR VGND sg13g2_nor3_2
X_3735_ net755 net505 _0602_ _0358_ VPWR VGND sg13g2_mux2_1
X_3666_ net771 _0551_ _1637_ VPWR VGND sg13g2_nor2_1
X_3597_ VGND VPWR net776 _1546_ _1571_ _0551_ sg13g2_a21oi_1
X_2617_ VGND VPWR _0896_ _0895_ _0595_ sg13g2_or2_1
X_2548_ _0745_ _0811_ _0740_ _0839_ VPWR VGND sg13g2_nand3_1
X_2479_ _0752_ _0775_ _0751_ _0776_ VPWR VGND sg13g2_nand3_1
X_4218_ net642 VGND VPWR net330 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[54\]
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
X_4149_ net654 VGND VPWR net433 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[69\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_43_316 VPWR VGND sg13g2_decap_8
XFILLER_11_202 VPWR VGND sg13g2_fill_1
Xclkload0 clkload0/Y clknet_leaf_55_clk VPWR VGND sg13g2_inv_2
XFILLER_4_935 VPWR VGND sg13g2_decap_8
XFILLER_3_423 VPWR VGND sg13g2_decap_4
XFILLER_47_644 VPWR VGND sg13g2_fill_2
XFILLER_46_121 VPWR VGND sg13g2_decap_8
XFILLER_46_165 VPWR VGND sg13g2_fill_1
XFILLER_28_891 VPWR VGND sg13g2_fill_2
XFILLER_43_894 VPWR VGND sg13g2_decap_8
XFILLER_30_588 VPWR VGND sg13g2_decap_4
XFILLER_7_740 VPWR VGND sg13g2_decap_8
X_3520_ _1495_ VPWR _1496_ VGND net799 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[32\]
+ sg13g2_o21ai_1
Xhold707 _0257_ VPWR VGND net1025 sg13g2_dlygate4sd3_1
Xhold718 u_usb_cdc.rstn VPWR VGND net1036 sg13g2_dlygate4sd3_1
Xhold729 _0259_ VPWR VGND net1047 sg13g2_dlygate4sd3_1
X_3451_ _1454_ net250 net580 VPWR VGND sg13g2_nand2_1
X_2402_ net755 u_usb_cdc.sie_out_data\[2\] _0702_ VPWR VGND sg13g2_nor2_2
X_3382_ net761 _1408_ _1409_ VPWR VGND sg13g2_nor2_1
XFILLER_3_990 VPWR VGND sg13g2_decap_8
X_2333_ _0634_ _0632_ _0633_ VPWR VGND sg13g2_nand2_1
X_2264_ _0566_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[1\] net794
+ VPWR VGND sg13g2_xnor2_1
XFILLER_38_600 VPWR VGND sg13g2_decap_8
X_2195_ VPWR _0497_ _0496_ VGND sg13g2_inv_1
XFILLER_26_806 VPWR VGND sg13g2_fill_1
X_4003_ _1881_ VPWR _0435_ VGND _1876_ _1882_ sg13g2_o21ai_1
XFILLER_26_817 VPWR VGND sg13g2_decap_8
XFILLER_34_872 VPWR VGND sg13g2_fill_1
XFILLER_34_894 VPWR VGND sg13g2_fill_1
X_3718_ net590 _1683_ net764 _1685_ VPWR VGND sg13g2_nand3_1
X_3649_ _1621_ _1620_ _1544_ _1619_ _1618_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_437 VPWR VGND sg13g2_decap_8
Xhold12 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[6\] VPWR VGND
+ net54 sg13g2_dlygate4sd3_1
Xhold23 _0211_ VPWR VGND net65 sg13g2_dlygate4sd3_1
XFILLER_29_23 VPWR VGND sg13g2_fill_2
Xhold45 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[54\] VPWR VGND
+ net87 sg13g2_dlygate4sd3_1
Xhold34 _0092_ VPWR VGND net76 sg13g2_dlygate4sd3_1
Xhold56 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[37\] VPWR VGND
+ net98 sg13g2_dlygate4sd3_1
Xhold89 _0127_ VPWR VGND net131 sg13g2_dlygate4sd3_1
Xhold78 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[66\] VPWR VGND
+ net120 sg13g2_dlygate4sd3_1
Xhold67 _0212_ VPWR VGND net109 sg13g2_dlygate4sd3_1
XFILLER_45_22 VPWR VGND sg13g2_fill_1
XFILLER_45_11 VPWR VGND sg13g2_fill_1
XFILLER_28_154 VPWR VGND sg13g2_decap_8
XFILLER_44_625 VPWR VGND sg13g2_fill_2
XFILLER_25_883 VPWR VGND sg13g2_decap_4
XFILLER_12_544 VPWR VGND sg13g2_fill_1
XFILLER_40_886 VPWR VGND sg13g2_decap_8
XFILLER_8_548 VPWR VGND sg13g2_decap_4
XFILLER_4_732 VPWR VGND sg13g2_decap_8
XFILLER_3_220 VPWR VGND sg13g2_decap_4
XFILLER_3_253 VPWR VGND sg13g2_fill_1
XFILLER_3_286 VPWR VGND sg13g2_decap_8
XFILLER_48_931 VPWR VGND sg13g2_decap_8
XFILLER_35_658 VPWR VGND sg13g2_fill_1
XFILLER_22_308 VPWR VGND sg13g2_decap_8
XFILLER_31_820 VPWR VGND sg13g2_fill_1
X_2951_ _1120_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ net603 VPWR VGND sg13g2_nand2_1
XFILLER_15_382 VPWR VGND sg13g2_fill_2
XFILLER_31_831 VPWR VGND sg13g2_decap_8
X_2882_ _1093_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ _1082_ VPWR VGND sg13g2_nand2_1
XFILLER_30_385 VPWR VGND sg13g2_fill_2
X_3503_ _0332_ net572 _0517_ net575 _1944_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_581 VPWR VGND sg13g2_fill_2
Xhold504 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[17\] VPWR
+ VGND net546 sg13g2_dlygate4sd3_1
Xhold526 _0362_ VPWR VGND net844 sg13g2_dlygate4sd3_1
Xhold515 _0955_ VPWR VGND net557 sg13g2_dlygate4sd3_1
Xhold559 _0249_ VPWR VGND net877 sg13g2_dlygate4sd3_1
Xhold537 _0293_ VPWR VGND net855 sg13g2_dlygate4sd3_1
X_3434_ net942 _0869_ _1446_ VPWR VGND sg13g2_nor2_1
Xhold548 u_usb_cdc.u_ctrl_endp.state_q\[5\] VPWR VGND net866 sg13g2_dlygate4sd3_1
XFILLER_44_1004 VPWR VGND sg13g2_decap_8
X_3365_ net415 _0711_ _1397_ _0282_ VPWR VGND sg13g2_mux2_1
X_3296_ _1274_ net819 net810 _1355_ VPWR VGND sg13g2_a21o_1
X_2316_ VPWR _0617_ _0616_ VGND sg13g2_inv_1
X_2247_ _0549_ net786 net785 VPWR VGND sg13g2_nand2_2
XFILLER_39_931 VPWR VGND sg13g2_decap_8
XFILLER_38_441 VPWR VGND sg13g2_decap_4
X_2178_ _0480_ net721 net757 VPWR VGND sg13g2_nand2_2
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_21_396 VPWR VGND sg13g2_fill_1
Xoutput24 net24 uio_out[2] VPWR VGND sg13g2_buf_1
Xoutput35 net35 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_757 VPWR VGND sg13g2_decap_8
XFILLER_49_739 VPWR VGND sg13g2_decap_8
XFILLER_0_256 VPWR VGND sg13g2_decap_8
XFILLER_45_912 VPWR VGND sg13g2_decap_8
XFILLER_17_625 VPWR VGND sg13g2_fill_2
XFILLER_45_989 VPWR VGND sg13g2_decap_8
XFILLER_44_477 VPWR VGND sg13g2_fill_1
XFILLER_32_628 VPWR VGND sg13g2_fill_2
XFILLER_40_650 VPWR VGND sg13g2_fill_1
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
X_3150_ _1232_ VPWR _0232_ VGND _1170_ _1229_ sg13g2_o21ai_1
X_3081_ _1195_ VPWR _0200_ VGND net720 net606 sg13g2_o21ai_1
X_2101_ VPWR _1979_ net180 VGND sg13g2_inv_1
XFILLER_11_4 VPWR VGND sg13g2_decap_8
X_2032_ VPWR _1911_ net829 VGND sg13g2_inv_1
XFILLER_35_433 VPWR VGND sg13g2_fill_2
XFILLER_36_989 VPWR VGND sg13g2_decap_8
X_3983_ VGND VPWR net210 net623 _0429_ _1868_ sg13g2_a21oi_1
X_2934_ _1114_ VPWR _0134_ VGND net707 _1089_ sg13g2_o21ai_1
XFILLER_31_650 VPWR VGND sg13g2_fill_1
X_2865_ _1081_ net162 _1080_ VPWR VGND sg13g2_nand2_1
Xhold301 _0950_ VPWR VGND net343 sg13g2_dlygate4sd3_1
X_2796_ _1032_ VPWR _0073_ VGND _1036_ _1037_ sg13g2_o21ai_1
Xhold334 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[39\] VPWR VGND
+ net376 sg13g2_dlygate4sd3_1
Xhold323 _0281_ VPWR VGND net365 sg13g2_dlygate4sd3_1
Xhold312 u_usb_cdc.u_sie.in_toggle_q\[2\] VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold367 u_usb_cdc.u_sie.crc16_q\[0\] VPWR VGND net409 sg13g2_dlygate4sd3_1
Xhold345 _1802_ VPWR VGND net387 sg13g2_dlygate4sd3_1
Xhold378 net15 VPWR VGND net420 sg13g2_dlygate4sd3_1
Xhold356 _0087_ VPWR VGND net398 sg13g2_dlygate4sd3_1
Xfanout825 net826 net825 VPWR VGND sg13g2_buf_1
Xfanout803 net804 net803 VPWR VGND sg13g2_buf_8
Xfanout814 net819 net814 VPWR VGND sg13g2_buf_8
X_4397_ net727 VGND VPWR _0399_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_2
X_3417_ net778 _0548_ net783 _1434_ VPWR VGND sg13g2_nand3_1
Xhold389 _0148_ VPWR VGND net431 sg13g2_dlygate4sd3_1
X_3348_ _0723_ _1387_ _1388_ VPWR VGND sg13g2_and2_1
Xfanout836 net837 net836 VPWR VGND sg13g2_buf_8
X_3279_ net818 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[39\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[47\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[55\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[63\] net811 _1344_
+ VPWR VGND sg13g2_mux4_1
XFILLER_41_403 VPWR VGND sg13g2_decap_4
XFILLER_26_477 VPWR VGND sg13g2_fill_1
XFILLER_6_849 VPWR VGND sg13g2_decap_8
XFILLER_1_554 VPWR VGND sg13g2_decap_8
XFILLER_49_547 VPWR VGND sg13g2_decap_8
XFILLER_17_444 VPWR VGND sg13g2_decap_8
XFILLER_45_797 VPWR VGND sg13g2_decap_8
XFILLER_32_403 VPWR VGND sg13g2_fill_2
XFILLER_33_915 VPWR VGND sg13g2_fill_1
XFILLER_17_499 VPWR VGND sg13g2_decap_8
XFILLER_9_643 VPWR VGND sg13g2_fill_1
XFILLER_13_694 VPWR VGND sg13g2_decap_8
XFILLER_9_665 VPWR VGND sg13g2_fill_2
X_2650_ VGND VPWR _2012_ _0920_ _0921_ _0442_ sg13g2_a21oi_1
X_2581_ _0864_ VPWR _0016_ VGND _1920_ _0863_ sg13g2_o21ai_1
X_4320_ net684 VGND VPWR net340 u_usb_cdc.u_sie.in_byte_q\[3\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_4251_ net649 VGND VPWR net961 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[3\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_2
X_3202_ _0966_ _0967_ _1274_ VPWR VGND sg13g2_nor2b_2
X_4182_ net645 VGND VPWR net322 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[18\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3133_ _1223_ net175 net627 VPWR VGND sg13g2_nand2_1
X_3064_ _1186_ VPWR _0192_ VGND net720 net608 sg13g2_o21ai_1
X_2015_ net761 _1894_ VPWR VGND sg13g2_inv_4
XFILLER_36_731 VPWR VGND sg13g2_decap_4
XFILLER_36_753 VPWR VGND sg13g2_decap_8
XFILLER_36_764 VPWR VGND sg13g2_fill_1
X_3966_ VPWR VGND _1854_ _1818_ _1808_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] _1855_
+ _0585_ sg13g2_a221oi_1
X_2917_ _1105_ VPWR _0126_ VGND _1070_ net615 sg13g2_o21ai_1
XFILLER_32_992 VPWR VGND sg13g2_decap_8
X_3897_ net386 net703 _1802_ VPWR VGND sg13g2_nor2_1
X_2848_ _1069_ net137 _1059_ VPWR VGND sg13g2_nand2_1
XFILLER_12_59 VPWR VGND sg13g2_decap_4
XFILLER_3_808 VPWR VGND sg13g2_decap_8
X_2779_ VGND VPWR _1022_ _1023_ _0070_ net924 sg13g2_a21oi_1
Xhold142 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[19\] VPWR VGND
+ net184 sg13g2_dlygate4sd3_1
Xhold153 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[43\] VPWR
+ VGND net195 sg13g2_dlygate4sd3_1
Xhold131 _0387_ VPWR VGND net173 sg13g2_dlygate4sd3_1
Xhold120 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[16\] VPWR VGND
+ net162 sg13g2_dlygate4sd3_1
Xhold164 u_usb_cdc.u_ctrl_endp.req_q\[10\] VPWR VGND net206 sg13g2_dlygate4sd3_1
Xhold175 _0176_ VPWR VGND net217 sg13g2_dlygate4sd3_1
Xhold186 _0191_ VPWR VGND net228 sg13g2_dlygate4sd3_1
X_4449_ net1 VGND VPWR net42 u_usb_cdc.rstn_sq\[1\] clknet_leaf_14_clk sg13g2_dfrbpq_1
Xfanout622 _1999_ net622 VPWR VGND sg13g2_buf_8
Xhold197 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[25\] VPWR
+ VGND net239 sg13g2_dlygate4sd3_1
Xfanout611 _1166_ net611 VPWR VGND sg13g2_buf_8
Xfanout600 _1739_ net600 VPWR VGND sg13g2_buf_8
Xfanout633 _0575_ net633 VPWR VGND sg13g2_buf_8
Xfanout655 net656 net655 VPWR VGND sg13g2_buf_8
Xfanout644 net645 net644 VPWR VGND sg13g2_buf_8
Xfanout666 net667 net666 VPWR VGND sg13g2_buf_8
Xfanout688 net689 net688 VPWR VGND sg13g2_buf_8
Xfanout677 net678 net677 VPWR VGND sg13g2_buf_8
Xfanout699 net700 net699 VPWR VGND sg13g2_buf_8
XFILLER_2_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_89 VPWR VGND sg13g2_decap_8
XFILLER_26_296 VPWR VGND sg13g2_decap_4
XFILLER_5_145 VPWR VGND sg13g2_decap_4
XFILLER_2_830 VPWR VGND sg13g2_decap_8
XFILLER_1_351 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_18_720 VPWR VGND sg13g2_decap_4
X_3820_ _1748_ _1750_ _0384_ VPWR VGND sg13g2_and2_1
X_3751_ net957 _1698_ _1695_ _0367_ VPWR VGND sg13g2_mux2_1
X_2702_ net51 net48 _0041_ VPWR VGND sg13g2_and2_1
X_3682_ _1912_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[46\] _1652_
+ VPWR VGND sg13g2_nor2_1
X_2633_ _0906_ VPWR _0028_ VGND _1957_ _0872_ sg13g2_o21ai_1
X_2564_ _0638_ _0681_ _1928_ _0853_ VPWR VGND _0851_ sg13g2_nand4_1
X_4303_ net691 VGND VPWR _0305_ u_usb_cdc.endp\[2\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_2495_ _0730_ VPWR _0792_ VGND _0479_ _0788_ sg13g2_o21ai_1
X_4234_ net639 VGND VPWR net117 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[70\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4165_ net661 VGND VPWR _0168_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[1\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3116_ net276 net604 _1214_ VPWR VGND sg13g2_nor2_1
X_4096_ net651 VGND VPWR net163 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[16\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3047_ net299 net612 _1175_ VPWR VGND sg13g2_nor2_1
XFILLER_23_288 VPWR VGND sg13g2_decap_4
X_3949_ net702 _1839_ _1840_ VPWR VGND sg13g2_nor2_1
XFILLER_24_1024 VPWR VGND sg13g2_decap_4
XFILLER_46_358 VPWR VGND sg13g2_fill_2
XFILLER_9_49 VPWR VGND sg13g2_fill_1
XFILLER_14_288 VPWR VGND sg13g2_fill_1
XFILLER_30_726 VPWR VGND sg13g2_fill_2
XFILLER_11_973 VPWR VGND sg13g2_decap_8
XFILLER_31_1017 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_955 VPWR VGND sg13g2_decap_8
X_2280_ u_usb_cdc.u_sie.phy_state_q\[2\] net186 u_usb_cdc.u_sie.phy_state_q\[3\] _0582_
+ VPWR VGND sg13g2_nor3_1
XFILLER_37_314 VPWR VGND sg13g2_decap_8
XFILLER_45_391 VPWR VGND sg13g2_fill_2
X_3803_ _1961_ _1980_ _1737_ VPWR VGND sg13g2_nor2_1
XFILLER_33_597 VPWR VGND sg13g2_decap_4
X_3734_ net756 net374 net589 _0357_ VPWR VGND sg13g2_mux2_1
X_3665_ _1918_ _0541_ _0670_ _1636_ VPWR VGND sg13g2_nor3_1
X_2616_ _0895_ _1990_ _0578_ VPWR VGND sg13g2_nand2_1
X_3596_ VGND VPWR net716 _1510_ _1570_ _1569_ sg13g2_a21oi_1
XFILLER_47_1024 VPWR VGND sg13g2_fill_1
XFILLER_0_619 VPWR VGND sg13g2_decap_8
X_2547_ _0838_ net206 _0692_ VPWR VGND sg13g2_nand2_1
X_2478_ u_usb_cdc.u_ctrl_endp.req_q\[3\] u_usb_cdc.u_ctrl_endp.req_q\[10\] u_usb_cdc.u_ctrl_endp.req_q\[9\]
+ _0775_ VPWR VGND sg13g2_nor3_1
X_4217_ net642 VGND VPWR net501 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[53\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_29_815 VPWR VGND sg13g2_decap_4
X_4148_ net668 VGND VPWR net449 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[68\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_44_829 VPWR VGND sg13g2_decap_8
XFILLER_28_358 VPWR VGND sg13g2_fill_2
X_4079_ net650 VGND VPWR _0082_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_24_531 VPWR VGND sg13g2_decap_8
XFILLER_12_748 VPWR VGND sg13g2_fill_2
Xclkload1 clknet_leaf_48_clk clkload1/Y VPWR VGND sg13g2_inv_4
XFILLER_20_792 VPWR VGND sg13g2_decap_8
XFILLER_4_914 VPWR VGND sg13g2_decap_8
XFILLER_3_402 VPWR VGND sg13g2_decap_8
XFILLER_46_111 VPWR VGND sg13g2_fill_1
XFILLER_15_520 VPWR VGND sg13g2_fill_1
XFILLER_34_339 VPWR VGND sg13g2_fill_2
XFILLER_15_531 VPWR VGND sg13g2_fill_1
XFILLER_43_873 VPWR VGND sg13g2_decap_8
XFILLER_11_792 VPWR VGND sg13g2_fill_2
Xhold719 u_usb_cdc.u_ctrl_endp.state_q\[2\] VPWR VGND net1037 sg13g2_dlygate4sd3_1
Xhold708 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[1\] VPWR VGND
+ net1026 sg13g2_dlygate4sd3_1
X_3450_ _1453_ VPWR _0311_ VGND _1898_ net581 sg13g2_o21ai_1
XFILLER_7_796 VPWR VGND sg13g2_decap_8
X_3381_ _0673_ VPWR _1408_ VGND _1900_ _0752_ sg13g2_o21ai_1
X_2401_ net841 u_usb_cdc.u_ctrl_endp.state_q\[6\] _0557_ _0681_ _0701_ VPWR VGND sg13g2_or4_1
X_2332_ _0633_ u_usb_cdc.u_ctrl_endp.state_q\[7\] _0605_ VPWR VGND sg13g2_nand2_1
XFILLER_2_490 VPWR VGND sg13g2_fill_2
X_2263_ _0565_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[2\] net790
+ VPWR VGND sg13g2_xnor2_1
XFILLER_38_612 VPWR VGND sg13g2_fill_2
X_4002_ _1879_ net333 _1882_ VPWR VGND sg13g2_xor2_1
X_2194_ _1925_ _0467_ u_usb_cdc.u_sie.pid_q\[2\] _0496_ VPWR VGND sg13g2_nand3_1
XFILLER_34_840 VPWR VGND sg13g2_fill_1
XFILLER_14_1023 VPWR VGND sg13g2_decap_4
XFILLER_21_567 VPWR VGND sg13g2_fill_2
X_3717_ _1684_ VPWR _0347_ VGND _1894_ net598 sg13g2_o21ai_1
X_3648_ _1525_ _1543_ _1620_ VPWR VGND sg13g2_and2_1
X_3579_ net777 _0550_ _0660_ _1554_ VPWR VGND sg13g2_nor3_1
XFILLER_0_416 VPWR VGND sg13g2_decap_8
XFILLER_1_939 VPWR VGND sg13g2_decap_8
Xhold13 _0173_ VPWR VGND net55 sg13g2_dlygate4sd3_1
XFILLER_29_35 VPWR VGND sg13g2_decap_4
Xhold46 _0137_ VPWR VGND net88 sg13g2_dlygate4sd3_1
Xhold35 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[35\] VPWR VGND
+ net77 sg13g2_dlygate4sd3_1
Xhold24 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[26\] VPWR VGND
+ net66 sg13g2_dlygate4sd3_1
Xhold68 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[42\] VPWR VGND
+ net110 sg13g2_dlygate4sd3_1
Xhold79 _0233_ VPWR VGND net121 sg13g2_dlygate4sd3_1
Xhold57 _0204_ VPWR VGND net99 sg13g2_dlygate4sd3_1
XFILLER_29_656 VPWR VGND sg13g2_fill_2
XFILLER_17_807 VPWR VGND sg13g2_fill_2
XFILLER_28_177 VPWR VGND sg13g2_fill_1
XFILLER_25_862 VPWR VGND sg13g2_decap_8
XFILLER_12_589 VPWR VGND sg13g2_fill_2
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_4_788 VPWR VGND sg13g2_decap_8
XFILLER_48_910 VPWR VGND sg13g2_decap_8
XFILLER_0_983 VPWR VGND sg13g2_decap_8
XFILLER_47_431 VPWR VGND sg13g2_fill_2
XFILLER_13_8 VPWR VGND sg13g2_fill_1
XFILLER_48_987 VPWR VGND sg13g2_decap_8
XFILLER_35_604 VPWR VGND sg13g2_fill_2
X_2950_ net462 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net603 _0145_ VPWR VGND sg13g2_mux2_1
XFILLER_16_884 VPWR VGND sg13g2_fill_1
X_2881_ _1092_ net93 _1080_ VPWR VGND sg13g2_nand2_1
XFILLER_42_180 VPWR VGND sg13g2_fill_2
XFILLER_30_331 VPWR VGND sg13g2_fill_2
XFILLER_31_876 VPWR VGND sg13g2_fill_1
XFILLER_31_887 VPWR VGND sg13g2_fill_1
X_3502_ _0331_ net573 _0516_ net577 _1945_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_593 VPWR VGND sg13g2_fill_1
Xhold505 _0184_ VPWR VGND net547 sg13g2_dlygate4sd3_1
Xhold527 u_usb_cdc.u_ctrl_endp.req_q\[8\] VPWR VGND net845 sg13g2_dlygate4sd3_1
Xhold516 _0036_ VPWR VGND net558 sg13g2_dlygate4sd3_1
Xhold538 u_usb_cdc.u_ctrl_endp.max_length_q\[1\] VPWR VGND net856 sg13g2_dlygate4sd3_1
Xhold549 _0015_ VPWR VGND net867 sg13g2_dlygate4sd3_1
X_3433_ net578 _1445_ _0302_ VPWR VGND sg13g2_and2_1
X_3364_ _0723_ _1396_ _1397_ VPWR VGND sg13g2_and2_1
X_3295_ net810 _1274_ net819 _1354_ VPWR VGND sg13g2_nand3_1
X_2315_ _0616_ _0571_ _0615_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_910 VPWR VGND sg13g2_decap_8
X_2246_ _1915_ net715 _0548_ VPWR VGND sg13g2_nor2_2
XFILLER_38_464 VPWR VGND sg13g2_decap_8
XFILLER_39_987 VPWR VGND sg13g2_decap_8
X_2177_ net760 net757 _0479_ VPWR VGND sg13g2_nor2_1
XFILLER_26_615 VPWR VGND sg13g2_decap_8
XFILLER_25_125 VPWR VGND sg13g2_decap_8
XFILLER_25_147 VPWR VGND sg13g2_decap_8
XFILLER_41_629 VPWR VGND sg13g2_decap_8
XFILLER_22_832 VPWR VGND sg13g2_decap_8
XFILLER_21_375 VPWR VGND sg13g2_decap_8
Xoutput25 net25 uio_out[3] VPWR VGND sg13g2_buf_1
Xoutput14 net14 uio_oe[0] VPWR VGND sg13g2_buf_1
Xoutput36 net36 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_736 VPWR VGND sg13g2_decap_8
XFILLER_0_213 VPWR VGND sg13g2_fill_2
XFILLER_49_718 VPWR VGND sg13g2_decap_8
XFILLER_29_420 VPWR VGND sg13g2_decap_4
XFILLER_44_423 VPWR VGND sg13g2_fill_1
XFILLER_45_968 VPWR VGND sg13g2_decap_8
XFILLER_44_434 VPWR VGND sg13g2_decap_4
XFILLER_8_346 VPWR VGND sg13g2_decap_8
XFILLER_12_375 VPWR VGND sg13g2_fill_2
X_2100_ VPWR _1978_ net102 VGND sg13g2_inv_1
XFILLER_0_780 VPWR VGND sg13g2_decap_8
X_3080_ _1195_ net188 net606 VPWR VGND sg13g2_nand2_1
X_2031_ _1910_ net835 VPWR VGND sg13g2_inv_2
XFILLER_48_784 VPWR VGND sg13g2_decap_8
XFILLER_47_250 VPWR VGND sg13g2_fill_2
XFILLER_36_968 VPWR VGND sg13g2_decap_8
X_3982_ net210 _1824_ _1868_ VPWR VGND sg13g2_nor2_1
X_2933_ _1114_ net159 _1110_ VPWR VGND sg13g2_nand2_1
XFILLER_44_990 VPWR VGND sg13g2_decap_8
X_2864_ _1080_ _1079_ VPWR VGND net616 sg13g2_nand2b_2
X_2795_ _1037_ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] net623 net743 _1893_ VPWR VGND
+ sg13g2_a22oi_1
XFILLER_11_1015 VPWR VGND sg13g2_decap_8
Xhold302 _0033_ VPWR VGND net344 sg13g2_dlygate4sd3_1
Xhold335 _0122_ VPWR VGND net377 sg13g2_dlygate4sd3_1
Xhold324 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[13\] VPWR VGND net366 sg13g2_dlygate4sd3_1
Xhold313 _1025_ VPWR VGND net355 sg13g2_dlygate4sd3_1
Xhold368 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[29\] VPWR VGND
+ net410 sg13g2_dlygate4sd3_1
Xhold357 u_usb_cdc.sie_out_data\[0\] VPWR VGND net399 sg13g2_dlygate4sd3_1
Xhold346 _0410_ VPWR VGND net388 sg13g2_dlygate4sd3_1
Xfanout804 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[0\] net804
+ VPWR VGND sg13g2_buf_8
Xfanout815 net816 net815 VPWR VGND sg13g2_buf_8
X_4396_ net725 VGND VPWR net190 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[17\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xhold379 _0356_ VPWR VGND net421 sg13g2_dlygate4sd3_1
X_3416_ _1433_ net778 _1424_ VPWR VGND sg13g2_nand2_1
Xfanout826 net1065 net826 VPWR VGND sg13g2_buf_8
X_3347_ _1386_ VPWR _1387_ VGND net751 _0778_ sg13g2_o21ai_1
Xfanout837 u_usb_cdc.u_sie.phy_state_q\[6\] net837 VPWR VGND sg13g2_buf_8
X_3278_ _0249_ _1343_ _1342_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_902 VPWR VGND sg13g2_fill_2
XFILLER_39_762 VPWR VGND sg13g2_fill_1
XFILLER_26_412 VPWR VGND sg13g2_decap_8
X_2229_ VGND VPWR _0499_ _0530_ _0531_ net746 sg13g2_a21oi_1
XFILLER_26_434 VPWR VGND sg13g2_fill_1
XFILLER_42_949 VPWR VGND sg13g2_decap_8
XFILLER_10_835 VPWR VGND sg13g2_fill_1
XFILLER_21_161 VPWR VGND sg13g2_fill_1
XFILLER_6_828 VPWR VGND sg13g2_decap_8
XFILLER_1_533 VPWR VGND sg13g2_decap_8
XFILLER_49_526 VPWR VGND sg13g2_decap_8
XFILLER_29_272 VPWR VGND sg13g2_fill_2
XFILLER_45_743 VPWR VGND sg13g2_decap_8
XFILLER_17_423 VPWR VGND sg13g2_fill_2
XFILLER_18_979 VPWR VGND sg13g2_decap_4
XFILLER_29_294 VPWR VGND sg13g2_fill_1
XFILLER_45_776 VPWR VGND sg13g2_decap_8
XFILLER_17_478 VPWR VGND sg13g2_decap_4
XFILLER_32_448 VPWR VGND sg13g2_decap_4
XFILLER_9_600 VPWR VGND sg13g2_fill_1
XFILLER_13_662 VPWR VGND sg13g2_fill_1
XFILLER_34_1015 VPWR VGND sg13g2_decap_8
XFILLER_41_982 VPWR VGND sg13g2_decap_8
XFILLER_13_684 VPWR VGND sg13g2_fill_2
X_2580_ _0638_ _0681_ net993 _0864_ VPWR VGND _0851_ sg13g2_nand4_1
XFILLER_5_883 VPWR VGND sg13g2_decap_8
X_4250_ net654 VGND VPWR net984 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[2\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_2
X_4181_ net645 VGND VPWR net547 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[17\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
X_3201_ net578 net1017 _1273_ _0242_ VPWR VGND sg13g2_a21o_1
X_3132_ _1222_ VPWR _0224_ VGND net720 net627 sg13g2_o21ai_1
X_3063_ _1186_ net239 net608 VPWR VGND sg13g2_nand2_1
X_2014_ VPWR _1893_ net308 VGND sg13g2_inv_1
XFILLER_36_798 VPWR VGND sg13g2_fill_2
XFILLER_23_448 VPWR VGND sg13g2_decap_8
X_3965_ _1854_ _1852_ _1853_ VPWR VGND sg13g2_nand2_1
XFILLER_23_459 VPWR VGND sg13g2_fill_1
X_2916_ _1105_ net149 _1101_ VPWR VGND sg13g2_nand2_1
X_3896_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] net852 _0448_ _0409_ VPWR VGND sg13g2_mux2_1
XFILLER_32_971 VPWR VGND sg13g2_decap_8
X_2847_ _1067_ VPWR _0093_ VGND net616 _1068_ sg13g2_o21ai_1
Xhold110 _0097_ VPWR VGND net152 sg13g2_dlygate4sd3_1
X_2778_ net739 _0990_ _1023_ VPWR VGND sg13g2_and2_1
Xhold143 _0102_ VPWR VGND net185 sg13g2_dlygate4sd3_1
Xhold132 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[34\] VPWR
+ VGND net174 sg13g2_dlygate4sd3_1
Xhold121 _0099_ VPWR VGND net163 sg13g2_dlygate4sd3_1
Xhold165 _0000_ VPWR VGND net207 sg13g2_dlygate4sd3_1
Xhold154 _0210_ VPWR VGND net196 sg13g2_dlygate4sd3_1
Xhold176 u_usb_cdc.u_sie.addr_q\[0\] VPWR VGND net218 sg13g2_dlygate4sd3_1
X_4448_ net1 VGND VPWR net45 u_usb_cdc.rstn clknet_leaf_14_clk sg13g2_dfrbpq_1
Xhold198 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[36\] VPWR
+ VGND net240 sg13g2_dlygate4sd3_1
Xfanout612 _1166_ net612 VPWR VGND sg13g2_buf_8
Xfanout601 _1275_ net601 VPWR VGND sg13g2_buf_8
Xhold187 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[7\] VPWR VGND
+ net229 sg13g2_dlygate4sd3_1
Xfanout623 _1998_ net623 VPWR VGND sg13g2_buf_8
Xfanout656 net657 net656 VPWR VGND sg13g2_buf_8
X_4379_ net723 VGND VPWR _0381_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[0\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_2
Xfanout645 net647 net645 VPWR VGND sg13g2_buf_8
Xfanout667 net701 net667 VPWR VGND sg13g2_buf_8
Xfanout634 _0572_ net634 VPWR VGND sg13g2_buf_8
Xfanout678 net690 net678 VPWR VGND sg13g2_buf_8
Xfanout689 net690 net689 VPWR VGND sg13g2_buf_8
XFILLER_15_927 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_fill_2
XFILLER_2_886 VPWR VGND sg13g2_decap_8
XFILLER_45_562 VPWR VGND sg13g2_fill_1
XFILLER_17_297 VPWR VGND sg13g2_fill_1
XFILLER_14_960 VPWR VGND sg13g2_decap_8
XFILLER_21_919 VPWR VGND sg13g2_fill_1
X_3750_ _1698_ _1003_ _1692_ VPWR VGND sg13g2_nand2_1
X_2701_ _0003_ _0959_ _0960_ VPWR VGND sg13g2_nand2_1
X_3681_ _1650_ VPWR _1651_ VGND net794 _1648_ sg13g2_o21ai_1
XFILLER_9_485 VPWR VGND sg13g2_fill_2
X_2632_ _0906_ net832 net595 VPWR VGND sg13g2_nand2_1
X_2563_ VPWR _0852_ _0851_ VGND sg13g2_inv_1
X_4302_ net681 VGND VPWR net959 u_usb_cdc.endp\[1\] clknet_leaf_36_clk sg13g2_dfrbpq_2
X_2494_ VGND VPWR _0791_ _0790_ _0729_ sg13g2_or2_1
X_4233_ net641 VGND VPWR net135 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[69\]
+ clknet_leaf_4_clk sg13g2_dfrbpq_1
X_4164_ net665 VGND VPWR net256 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[0\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_4095_ net669 VGND VPWR net92 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[15\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3115_ VGND VPWR _1170_ net604 _0216_ _1213_ sg13g2_a21oi_1
X_3046_ VGND VPWR net611 _1173_ _0186_ _1174_ sg13g2_a21oi_1
XFILLER_36_540 VPWR VGND sg13g2_decap_4
XFILLER_23_201 VPWR VGND sg13g2_fill_2
XFILLER_36_573 VPWR VGND sg13g2_fill_1
XFILLER_11_418 VPWR VGND sg13g2_fill_2
XFILLER_23_267 VPWR VGND sg13g2_decap_8
XFILLER_23_48 VPWR VGND sg13g2_decap_4
X_3948_ _1838_ VPWR _1839_ VGND u_usb_cdc.u_sie.u_phy_tx.data_q\[4\] _2002_ sg13g2_o21ai_1
X_3879_ VGND VPWR _1788_ _1789_ _1793_ net52 sg13g2_a21oi_1
XFILLER_2_105 VPWR VGND sg13g2_decap_4
XFILLER_24_1003 VPWR VGND sg13g2_decap_8
XFILLER_47_849 VPWR VGND sg13g2_decap_8
XFILLER_46_337 VPWR VGND sg13g2_fill_2
XFILLER_9_39 VPWR VGND sg13g2_fill_1
XFILLER_11_952 VPWR VGND sg13g2_decap_8
XFILLER_7_934 VPWR VGND sg13g2_decap_8
XFILLER_10_484 VPWR VGND sg13g2_fill_2
XFILLER_9_1008 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_8
XFILLER_49_142 VPWR VGND sg13g2_fill_2
XFILLER_46_893 VPWR VGND sg13g2_decap_8
X_3802_ _1734_ VPWR _0380_ VGND net516 _1736_ sg13g2_o21ai_1
XFILLER_14_790 VPWR VGND sg13g2_decap_4
X_3733_ net759 net420 net589 _0356_ VPWR VGND sg13g2_mux2_1
X_3664_ _1627_ VPWR _1635_ VGND net788 _1634_ sg13g2_o21ai_1
X_2615_ _0894_ net835 net592 VPWR VGND sg13g2_nand2_2
XFILLER_47_1003 VPWR VGND sg13g2_decap_8
X_3595_ VGND VPWR _0541_ _0549_ _1569_ net776 sg13g2_a21oi_1
X_2546_ _0836_ net949 _0837_ _0010_ VPWR VGND sg13g2_a21o_1
X_2477_ net736 VPWR _0774_ VGND _0761_ _0773_ sg13g2_o21ai_1
X_4216_ net660 VGND VPWR net324 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[52\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_4147_ net654 VGND VPWR net478 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[67\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_28_337 VPWR VGND sg13g2_fill_2
X_4078_ net650 VGND VPWR _0081_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_2
X_3029_ net823 _1150_ net752 _1163_ VPWR VGND sg13g2_nand3_1
XFILLER_37_882 VPWR VGND sg13g2_decap_4
Xclkload2 clknet_leaf_35_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_28_860 VPWR VGND sg13g2_fill_1
XFILLER_35_819 VPWR VGND sg13g2_fill_2
XFILLER_43_841 VPWR VGND sg13g2_decap_8
XFILLER_15_587 VPWR VGND sg13g2_fill_2
XFILLER_30_557 VPWR VGND sg13g2_decap_8
XFILLER_7_775 VPWR VGND sg13g2_decap_8
Xhold709 _1367_ VPWR VGND net1027 sg13g2_dlygate4sd3_1
X_2400_ _0700_ _0662_ net574 VPWR VGND sg13g2_nand2_1
X_3380_ net864 net568 _1407_ VPWR VGND sg13g2_nor2_1
X_2331_ net841 u_usb_cdc.u_ctrl_endp.state_q\[5\] u_usb_cdc.u_ctrl_endp.state_q\[6\]
+ _0632_ VPWR VGND sg13g2_nor3_1
X_2262_ _0564_ net803 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\]
+ VPWR VGND sg13g2_nand2b_1
X_4001_ _1881_ net333 net713 VPWR VGND sg13g2_nand2_1
X_2193_ _0495_ u_usb_cdc.u_sie.pid_q\[2\] _1925_ VPWR VGND sg13g2_nand2_1
XFILLER_38_657 VPWR VGND sg13g2_fill_1
XFILLER_33_373 VPWR VGND sg13g2_decap_8
XFILLER_14_1002 VPWR VGND sg13g2_decap_8
XFILLER_21_579 VPWR VGND sg13g2_fill_1
X_3716_ net590 _1683_ net766 _1684_ VPWR VGND sg13g2_nand3_1
X_3647_ _1619_ _0850_ _0552_ _0652_ _0544_ VPWR VGND sg13g2_a22oi_1
XFILLER_1_918 VPWR VGND sg13g2_decap_8
X_3578_ _1516_ _1548_ _1551_ _1552_ _1553_ VPWR VGND sg13g2_nor4_1
X_2529_ _0693_ _0767_ _0662_ _0824_ VPWR VGND sg13g2_nand3_1
Xhold14 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[45\] VPWR VGND
+ net56 sg13g2_dlygate4sd3_1
Xhold36 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[40\] VPWR VGND
+ net78 sg13g2_dlygate4sd3_1
Xhold47 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[17\] VPWR VGND
+ net89 sg13g2_dlygate4sd3_1
Xhold25 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[23\] VPWR VGND
+ net67 sg13g2_dlygate4sd3_1
Xhold69 _0125_ VPWR VGND net111 sg13g2_dlygate4sd3_1
Xhold58 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[68\] VPWR VGND
+ net100 sg13g2_dlygate4sd3_1
XFILLER_29_624 VPWR VGND sg13g2_decap_8
XFILLER_44_605 VPWR VGND sg13g2_fill_2
XFILLER_43_148 VPWR VGND sg13g2_fill_1
XFILLER_24_384 VPWR VGND sg13g2_fill_2
XFILLER_4_767 VPWR VGND sg13g2_decap_8
XFILLER_0_962 VPWR VGND sg13g2_decap_8
XFILLER_48_966 VPWR VGND sg13g2_decap_8
XFILLER_19_134 VPWR VGND sg13g2_fill_1
XFILLER_47_487 VPWR VGND sg13g2_decap_8
XFILLER_19_167 VPWR VGND sg13g2_fill_2
XFILLER_34_159 VPWR VGND sg13g2_fill_1
XFILLER_37_1024 VPWR VGND sg13g2_decap_4
XFILLER_15_384 VPWR VGND sg13g2_fill_1
X_2880_ _1090_ VPWR _0103_ VGND net824 _1091_ sg13g2_o21ai_1
XFILLER_30_354 VPWR VGND sg13g2_fill_1
XFILLER_30_365 VPWR VGND sg13g2_decap_8
XFILLER_30_387 VPWR VGND sg13g2_fill_1
Xhold506 u_usb_cdc.u_sie.crc16_q\[12\] VPWR VGND net548 sg13g2_dlygate4sd3_1
X_3501_ _0330_ _1484_ _0521_ net576 _1952_ VPWR VGND sg13g2_a22oi_1
XFILLER_7_583 VPWR VGND sg13g2_fill_1
Xhold517 net32 VPWR VGND net559 sg13g2_dlygate4sd3_1
Xhold539 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[2\] VPWR VGND
+ net857 sg13g2_dlygate4sd3_1
Xhold528 _0009_ VPWR VGND net846 sg13g2_dlygate4sd3_1
X_3432_ _1445_ _1239_ net769 VPWR VGND sg13g2_nand2b_1
X_3363_ _1386_ VPWR _1396_ VGND _0710_ _0784_ sg13g2_o21ai_1
X_3294_ VGND VPWR net814 _1274_ _0255_ _1353_ sg13g2_a21oi_1
X_2314_ _0573_ _0614_ _0615_ VPWR VGND sg13g2_nor2_1
X_2245_ _0547_ net787 VPWR VGND net782 sg13g2_nand2b_2
X_2176_ _0478_ net760 net757 VPWR VGND sg13g2_nand2_1
XFILLER_39_966 VPWR VGND sg13g2_decap_8
XFILLER_26_627 VPWR VGND sg13g2_decap_8
XFILLER_19_690 VPWR VGND sg13g2_fill_2
Xoutput15 net15 uio_oe[1] VPWR VGND sg13g2_buf_1
XFILLER_1_715 VPWR VGND sg13g2_decap_8
Xoutput26 net26 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput37 net37 usb_dn_en_o VPWR VGND sg13g2_buf_1
XFILLER_29_410 VPWR VGND sg13g2_decap_4
XFILLER_45_947 VPWR VGND sg13g2_decap_8
XFILLER_17_627 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_51_clk clknet_3_1__leaf_clk clknet_leaf_51_clk VPWR VGND sg13g2_buf_8
XFILLER_48_763 VPWR VGND sg13g2_decap_8
X_2030_ VPWR _1909_ net1034 VGND sg13g2_inv_1
XFILLER_36_947 VPWR VGND sg13g2_decap_8
X_3981_ net622 net368 _1867_ _0428_ VPWR VGND sg13g2_a21o_1
X_2932_ _1113_ VPWR _0133_ VGND net707 _1087_ sg13g2_o21ai_1
XFILLER_16_693 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_42_clk clknet_3_5__leaf_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
X_2863_ net828 net827 _1079_ VPWR VGND sg13g2_nor2b_2
XFILLER_30_195 VPWR VGND sg13g2_fill_1
X_2794_ VGND VPWR _2006_ _1035_ _1036_ _1996_ sg13g2_a21oi_1
XFILLER_7_61 VPWR VGND sg13g2_fill_2
Xhold325 _0394_ VPWR VGND net367 sg13g2_dlygate4sd3_1
Xhold303 u_usb_cdc.u_ctrl_endp.dev_state_q\[1\] VPWR VGND net345 sg13g2_dlygate4sd3_1
Xhold314 _0071_ VPWR VGND net356 sg13g2_dlygate4sd3_1
Xhold369 _0112_ VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold358 u_usb_cdc.u_sie.u_phy_tx.data_q\[6\] VPWR VGND net400 sg13g2_dlygate4sd3_1
Xhold347 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[16\] VPWR
+ VGND net389 sg13g2_dlygate4sd3_1
Xhold336 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[0\] VPWR VGND
+ net378 sg13g2_dlygate4sd3_1
Xfanout805 net806 net805 VPWR VGND sg13g2_buf_8
Xfanout816 net817 net816 VPWR VGND sg13g2_buf_8
X_4395_ net726 VGND VPWR _0397_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_2
X_3415_ _1431_ VPWR _0297_ VGND _1426_ _1432_ sg13g2_o21ai_1
Xfanout827 net1053 net827 VPWR VGND sg13g2_buf_8
X_3346_ _1386_ net738 net619 VPWR VGND sg13g2_nand2_1
Xfanout838 net939 net838 VPWR VGND sg13g2_buf_8
X_3277_ _1343_ _1296_ net116 net602 net876 VPWR VGND sg13g2_a22oi_1
X_2228_ VGND VPWR net833 _0529_ _0530_ net836 sg13g2_a21oi_1
X_2159_ u_usb_cdc.addr\[4\] net754 _0461_ VPWR VGND sg13g2_xor2_1
XFILLER_42_928 VPWR VGND sg13g2_decap_8
XFILLER_13_118 VPWR VGND sg13g2_fill_2
XFILLER_42_14 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_33_clk clknet_3_7__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
XFILLER_42_69 VPWR VGND sg13g2_fill_1
XFILLER_21_151 VPWR VGND sg13g2_fill_2
XFILLER_6_807 VPWR VGND sg13g2_decap_8
XFILLER_1_512 VPWR VGND sg13g2_decap_8
XFILLER_49_505 VPWR VGND sg13g2_decap_8
XFILLER_1_589 VPWR VGND sg13g2_decap_8
XFILLER_45_722 VPWR VGND sg13g2_decap_8
XFILLER_17_413 VPWR VGND sg13g2_decap_4
XFILLER_18_958 VPWR VGND sg13g2_decap_8
XFILLER_17_457 VPWR VGND sg13g2_fill_1
XFILLER_32_405 VPWR VGND sg13g2_fill_1
XFILLER_44_287 VPWR VGND sg13g2_fill_2
XFILLER_44_276 VPWR VGND sg13g2_decap_8
XFILLER_41_961 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_3_6__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_8_177 VPWR VGND sg13g2_fill_2
XFILLER_5_862 VPWR VGND sg13g2_decap_8
X_4180_ net645 VGND VPWR net390 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[16\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3200_ VGND VPWR _1269_ _1272_ _1273_ net578 sg13g2_a21oi_1
X_3131_ _1222_ net199 net627 VPWR VGND sg13g2_nand2_1
X_3062_ _1185_ VPWR _0191_ VGND net721 net608 sg13g2_o21ai_1
XFILLER_24_928 VPWR VGND sg13g2_fill_1
XFILLER_35_265 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_3_2__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
XFILLER_32_950 VPWR VGND sg13g2_decap_8
X_3964_ _1853_ u_usb_cdc.u_sie.data_q\[5\] net835 _1923_ net830 VPWR VGND sg13g2_a22oi_1
X_2915_ _1104_ VPWR _0125_ VGND _1068_ net615 sg13g2_o21ai_1
X_3895_ VGND VPWR _1935_ _0448_ _0408_ _1801_ sg13g2_a21oi_1
X_2846_ _1068_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2777_ _0993_ net479 net842 _1022_ VPWR VGND sg13g2_a21o_1
Xhold100 _0206_ VPWR VGND net142 sg13g2_dlygate4sd3_1
Xhold111 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[12\] VPWR
+ VGND net153 sg13g2_dlygate4sd3_1
Xhold122 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[59\] VPWR
+ VGND net164 sg13g2_dlygate4sd3_1
Xhold133 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[58\] VPWR
+ VGND net175 sg13g2_dlygate4sd3_1
Xhold144 u_usb_cdc.u_sie.phy_state_q\[5\] VPWR VGND net186 sg13g2_dlygate4sd3_1
X_4447_ net726 VGND VPWR _0040_ u_usb_cdc.clk_cnt_q\[1\] clknet_leaf_42_clk sg13g2_dfrbpq_1
Xhold155 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[46\] VPWR
+ VGND net197 sg13g2_dlygate4sd3_1
Xhold177 _1030_ VPWR VGND net219 sg13g2_dlygate4sd3_1
Xhold166 _0050_ VPWR VGND net208 sg13g2_dlygate4sd3_1
Xhold188 u_usb_cdc.u_sie.in_byte_q\[2\] VPWR VGND net230 sg13g2_dlygate4sd3_1
Xhold199 _0203_ VPWR VGND net241 sg13g2_dlygate4sd3_1
Xfanout613 net614 net613 VPWR VGND sg13g2_buf_8
Xfanout602 _1275_ net602 VPWR VGND sg13g2_buf_1
Xfanout624 net625 net624 VPWR VGND sg13g2_buf_8
Xfanout646 net647 net646 VPWR VGND sg13g2_buf_8
Xfanout635 _0450_ net635 VPWR VGND sg13g2_buf_8
X_4378_ net732 VGND VPWR net517 _0056_ clknet_leaf_32_clk sg13g2_dfrbpq_2
Xfanout657 net658 net657 VPWR VGND sg13g2_buf_8
X_3329_ VGND VPWR net720 _1377_ _0264_ _1379_ sg13g2_a21oi_1
Xfanout679 net682 net679 VPWR VGND sg13g2_buf_8
Xfanout668 net671 net668 VPWR VGND sg13g2_buf_8
XFILLER_15_906 VPWR VGND sg13g2_fill_1
XFILLER_10_644 VPWR VGND sg13g2_decap_8
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_49_313 VPWR VGND sg13g2_decap_8
XFILLER_1_386 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_32_224 VPWR VGND sg13g2_decap_4
XFILLER_33_758 VPWR VGND sg13g2_decap_8
X_2700_ _0713_ _0780_ _0695_ _0960_ VPWR VGND sg13g2_nand3_1
X_3680_ VGND VPWR net793 _1649_ _1650_ net789 sg13g2_a21oi_1
X_2631_ _0904_ VPWR _0027_ VGND _0872_ _0905_ sg13g2_o21ai_1
X_2562_ net953 _0649_ _0850_ _0851_ VPWR VGND sg13g2_nor3_1
X_4301_ net686 VGND VPWR net943 u_usb_cdc.endp\[0\] clknet_leaf_35_clk sg13g2_dfrbpq_2
X_2493_ VPWR VGND _0789_ _0731_ _0728_ net618 _0790_ _0727_ sg13g2_a221oi_1
X_4232_ net639 VGND VPWR net101 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[68\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_4_clk clknet_3_0__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ net673 VGND VPWR net336 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[3\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_2
X_4094_ net670 VGND VPWR net152 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[14\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3114_ net416 net604 _1213_ VPWR VGND sg13g2_nor2_1
X_3045_ net440 net611 _1174_ VPWR VGND sg13g2_nor2_1
XFILLER_12_909 VPWR VGND sg13g2_decap_8
XFILLER_17_1022 VPWR VGND sg13g2_decap_8
X_3947_ _1838_ _2004_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] VPWR VGND sg13g2_nand2b_1
X_3878_ _1791_ net295 _0400_ VPWR VGND sg13g2_nor2_1
X_2829_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net424 _1058_ _0085_ VPWR VGND sg13g2_mux2_1
XFILLER_3_8 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_fill_2
XFILLER_47_828 VPWR VGND sg13g2_decap_8
XFILLER_42_544 VPWR VGND sg13g2_decap_8
XFILLER_42_533 VPWR VGND sg13g2_fill_2
XFILLER_14_257 VPWR VGND sg13g2_decap_4
XFILLER_11_931 VPWR VGND sg13g2_decap_8
XFILLER_23_780 VPWR VGND sg13g2_fill_1
XFILLER_10_452 VPWR VGND sg13g2_fill_2
XFILLER_7_913 VPWR VGND sg13g2_decap_8
XFILLER_6_423 VPWR VGND sg13g2_decap_8
XFILLER_6_478 VPWR VGND sg13g2_fill_2
XFILLER_2_662 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_46_872 VPWR VGND sg13g2_decap_8
XFILLER_45_360 VPWR VGND sg13g2_decap_4
XFILLER_18_585 VPWR VGND sg13g2_decap_8
XFILLER_45_393 VPWR VGND sg13g2_fill_1
X_3801_ _1736_ _0443_ _0930_ VPWR VGND sg13g2_nand2_1
XFILLER_9_261 VPWR VGND sg13g2_decap_8
X_3732_ net761 net412 net589 _0355_ VPWR VGND sg13g2_mux2_1
X_3663_ _1633_ VPWR _1634_ VGND net789 _1628_ sg13g2_o21ai_1
XFILLER_9_283 VPWR VGND sg13g2_fill_1
X_2614_ net595 net525 _0893_ _0022_ VPWR VGND sg13g2_a21o_1
X_3594_ _1560_ VPWR _1568_ VGND net788 _1567_ sg13g2_o21ai_1
X_2545_ _0480_ _0728_ _0741_ _0788_ _0837_ VPWR VGND sg13g2_nor4_1
X_2476_ _0764_ _0765_ _0762_ _0773_ VPWR VGND _0772_ sg13g2_nand4_1
X_4215_ net639 VGND VPWR net326 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[51\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
X_4146_ net653 VGND VPWR net465 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[66\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4077_ net650 VGND VPWR _0080_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3028_ _1162_ net180 _1146_ VPWR VGND sg13g2_nand2_1
Xclkload3 clknet_leaf_29_clk clkload3/X VPWR VGND sg13g2_buf_8
XFILLER_20_761 VPWR VGND sg13g2_decap_8
XFILLER_4_949 VPWR VGND sg13g2_decap_8
XFILLER_3_459 VPWR VGND sg13g2_decap_8
XFILLER_3_437 VPWR VGND sg13g2_decap_4
XFILLER_42_363 VPWR VGND sg13g2_decap_4
XFILLER_11_794 VPWR VGND sg13g2_fill_1
XFILLER_7_754 VPWR VGND sg13g2_decap_8
X_2330_ VPWR VGND _0630_ _0573_ _0629_ _0620_ _0631_ _0621_ sg13g2_a221oi_1
XFILLER_2_492 VPWR VGND sg13g2_fill_1
X_2261_ VGND VPWR _0554_ _0561_ _0563_ _0562_ sg13g2_a21oi_1
XFILLER_27_4 VPWR VGND sg13g2_fill_2
X_4000_ _1878_ VPWR _0434_ VGND _1876_ _1880_ sg13g2_o21ai_1
X_2192_ _0477_ _0487_ _0491_ _0493_ _0494_ VPWR VGND sg13g2_and4_1
XFILLER_1_74 VPWR VGND sg13g2_fill_1
XFILLER_38_669 VPWR VGND sg13g2_decap_8
XFILLER_18_371 VPWR VGND sg13g2_decap_4
XFILLER_25_308 VPWR VGND sg13g2_fill_2
XFILLER_45_190 VPWR VGND sg13g2_fill_2
XFILLER_33_363 VPWR VGND sg13g2_decap_4
XFILLER_21_547 VPWR VGND sg13g2_decap_8
XFILLER_21_569 VPWR VGND sg13g2_fill_1
X_3715_ _1683_ _1957_ _0905_ VPWR VGND sg13g2_nand2_2
XFILLER_20_28 VPWR VGND sg13g2_fill_2
X_3646_ _1516_ _1617_ _1618_ VPWR VGND sg13g2_nor2_1
X_3577_ VPWR VGND _1430_ _1440_ _1510_ _0541_ _1552_ _1505_ sg13g2_a221oi_1
X_2528_ net574 net617 _0657_ _0823_ VPWR VGND sg13g2_nand3_1
Xhold15 _0128_ VPWR VGND net57 sg13g2_dlygate4sd3_1
Xhold37 _0207_ VPWR VGND net79 sg13g2_dlygate4sd3_1
X_2459_ VPWR _0756_ _0755_ VGND sg13g2_inv_1
Xhold26 _0106_ VPWR VGND net68 sg13g2_dlygate4sd3_1
Xhold59 _0235_ VPWR VGND net101 sg13g2_dlygate4sd3_1
Xhold48 _0100_ VPWR VGND net90 sg13g2_dlygate4sd3_1
X_4129_ net650 VGND VPWR net115 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[49\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_45_47 VPWR VGND sg13g2_fill_2
XFILLER_16_319 VPWR VGND sg13g2_decap_8
XFILLER_25_820 VPWR VGND sg13g2_decap_8
XFILLER_28_168 VPWR VGND sg13g2_decap_8
XFILLER_24_374 VPWR VGND sg13g2_fill_1
XFILLER_24_396 VPWR VGND sg13g2_fill_1
XFILLER_12_558 VPWR VGND sg13g2_decap_4
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_3_278 VPWR VGND sg13g2_fill_2
XFILLER_0_941 VPWR VGND sg13g2_decap_8
XFILLER_48_945 VPWR VGND sg13g2_decap_8
XFILLER_35_606 VPWR VGND sg13g2_fill_1
XFILLER_35_617 VPWR VGND sg13g2_fill_2
XFILLER_35_639 VPWR VGND sg13g2_fill_1
XFILLER_28_691 VPWR VGND sg13g2_fill_2
XFILLER_16_875 VPWR VGND sg13g2_decap_8
XFILLER_37_1003 VPWR VGND sg13g2_decap_8
XFILLER_30_300 VPWR VGND sg13g2_fill_1
XFILLER_30_333 VPWR VGND sg13g2_fill_1
X_3500_ _0329_ net573 _0506_ net576 _1953_ VPWR VGND sg13g2_a22oi_1
Xhold507 _0518_ VPWR VGND net549 sg13g2_dlygate4sd3_1
Xhold518 _0246_ VPWR VGND net560 sg13g2_dlygate4sd3_1
X_3431_ _1443_ VPWR _0301_ VGND _1426_ _1444_ sg13g2_o21ai_1
Xhold529 u_usb_cdc.u_sie.phy_state_q\[8\] VPWR VGND net847 sg13g2_dlygate4sd3_1
X_3362_ VGND VPWR _1901_ net571 _0281_ _1395_ sg13g2_a21oi_1
XFILLER_44_1018 VPWR VGND sg13g2_decap_8
X_2313_ u_usb_cdc.u_ctrl_endp.state_q\[2\] u_usb_cdc.u_ctrl_endp.state_q\[6\] _0557_
+ _0614_ VPWR VGND sg13g2_or3_1
X_3293_ VGND VPWR _1274_ _1286_ _1353_ net812 sg13g2_a21oi_1
X_2244_ net785 _0543_ _0544_ _0545_ _0546_ VPWR VGND sg13g2_and4_1
XFILLER_38_411 VPWR VGND sg13g2_fill_2
XFILLER_39_945 VPWR VGND sg13g2_decap_8
X_2175_ _0477_ u_usb_cdc.u_sie.data_q\[7\] _0476_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_190 VPWR VGND sg13g2_fill_2
XFILLER_21_333 VPWR VGND sg13g2_fill_2
XFILLER_21_355 VPWR VGND sg13g2_decap_8
XFILLER_31_16 VPWR VGND sg13g2_decap_4
X_3629_ VPWR VGND _1528_ _1489_ _1601_ net631 _1602_ _1591_ sg13g2_a221oi_1
Xoutput38 net38 usb_dn_tx_o VPWR VGND sg13g2_buf_1
Xoutput27 net27 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput16 net16 uio_oe[2] VPWR VGND sg13g2_buf_1
XFILLER_5_1023 VPWR VGND sg13g2_decap_4
XFILLER_45_926 VPWR VGND sg13g2_decap_8
XFILLER_25_661 VPWR VGND sg13g2_decap_4
XFILLER_13_812 VPWR VGND sg13g2_fill_1
XFILLER_13_834 VPWR VGND sg13g2_fill_2
XFILLER_12_322 VPWR VGND sg13g2_fill_2
XFILLER_12_377 VPWR VGND sg13g2_fill_1
XFILLER_48_742 VPWR VGND sg13g2_decap_8
XFILLER_47_285 VPWR VGND sg13g2_decap_4
X_3980_ VPWR VGND _1866_ _1825_ _1817_ net829 _1867_ net705 sg13g2_a221oi_1
X_2931_ _1113_ net124 _1110_ VPWR VGND sg13g2_nand2_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_2862_ _1077_ VPWR _0098_ VGND _1064_ _1078_ sg13g2_o21ai_1
XFILLER_31_664 VPWR VGND sg13g2_fill_1
XFILLER_30_174 VPWR VGND sg13g2_decap_8
X_2793_ VPWR VGND net702 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] _1994_ _1893_ _1035_
+ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] sg13g2_a221oi_1
XFILLER_8_882 VPWR VGND sg13g2_decap_8
XFILLER_7_73 VPWR VGND sg13g2_fill_1
XFILLER_7_84 VPWR VGND sg13g2_fill_2
Xhold304 u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\] VPWR VGND net346 sg13g2_dlygate4sd3_1
Xhold315 u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold326 _0057_ VPWR VGND net368 sg13g2_dlygate4sd3_1
Xhold359 _1862_ VPWR VGND net401 sg13g2_dlygate4sd3_1
Xhold348 _0183_ VPWR VGND net390 sg13g2_dlygate4sd3_1
X_3414_ _0549_ net783 _1432_ VPWR VGND sg13g2_xor2_1
Xhold337 _0083_ VPWR VGND net379 sg13g2_dlygate4sd3_1
X_4394_ net726 VGND VPWR _0396_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[15\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xfanout806 net1064 net806 VPWR VGND sg13g2_buf_8
Xfanout828 net1067 net828 VPWR VGND sg13g2_buf_8
X_3345_ net886 net364 _1384_ _0274_ VPWR VGND sg13g2_mux2_1
Xfanout817 net818 net817 VPWR VGND sg13g2_buf_8
Xfanout839 u_usb_cdc.u_sie.phy_state_q\[1\] net839 VPWR VGND sg13g2_buf_8
X_3276_ net805 net602 _1338_ _1341_ _1342_ VPWR VGND sg13g2_nor4_1
X_2227_ _0529_ net706 _0528_ VPWR VGND sg13g2_nand2_1
X_2158_ u_usb_cdc.addr\[1\] net758 _0460_ VPWR VGND sg13g2_xor2_1
XFILLER_26_425 VPWR VGND sg13g2_decap_8
XFILLER_42_907 VPWR VGND sg13g2_decap_8
X_2089_ VPWR _1967_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[40\]
+ VGND sg13g2_inv_1
XFILLER_35_992 VPWR VGND sg13g2_decap_8
XFILLER_21_130 VPWR VGND sg13g2_fill_2
XFILLER_21_141 VPWR VGND sg13g2_fill_2
XFILLER_1_568 VPWR VGND sg13g2_decap_8
XFILLER_27_1013 VPWR VGND sg13g2_decap_8
XFILLER_29_230 VPWR VGND sg13g2_decap_4
XFILLER_45_701 VPWR VGND sg13g2_decap_8
XFILLER_18_904 VPWR VGND sg13g2_fill_1
XFILLER_18_937 VPWR VGND sg13g2_decap_8
XFILLER_17_425 VPWR VGND sg13g2_fill_1
XFILLER_29_285 VPWR VGND sg13g2_decap_8
XFILLER_41_940 VPWR VGND sg13g2_decap_8
XFILLER_40_483 VPWR VGND sg13g2_decap_4
XFILLER_5_841 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_decap_4
X_3130_ _1221_ VPWR _0223_ VGND net721 net627 sg13g2_o21ai_1
X_3061_ _1185_ net227 net608 VPWR VGND sg13g2_nand2_1
X_3963_ _1852_ _1949_ net831 _1943_ net838 VPWR VGND sg13g2_a22oi_1
X_2914_ _1104_ net110 _1101_ VPWR VGND sg13g2_nand2_1
X_3894_ net913 _0448_ _1801_ VPWR VGND sg13g2_nor2_1
X_2845_ _1067_ net191 _1059_ VPWR VGND sg13g2_nand2_1
Xhold101 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[71\] VPWR
+ VGND net143 sg13g2_dlygate4sd3_1
X_2776_ _1021_ _1020_ _0574_ _1015_ net923 VPWR VGND sg13g2_a22oi_1
Xhold112 _0179_ VPWR VGND net154 sg13g2_dlygate4sd3_1
Xhold134 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[28\] VPWR
+ VGND net176 sg13g2_dlygate4sd3_1
Xhold123 u_usb_cdc.u_sie.in_zlp_q\[0\] VPWR VGND net165 sg13g2_dlygate4sd3_1
X_4446_ net726 VGND VPWR _0039_ u_usb_cdc.clk_cnt_q\[0\] clknet_leaf_42_clk sg13g2_dfrbpq_1
Xhold156 _0213_ VPWR VGND net198 sg13g2_dlygate4sd3_1
Xhold145 _0024_ VPWR VGND net187 sg13g2_dlygate4sd3_1
Xhold167 _0025_ VPWR VGND net209 sg13g2_dlygate4sd3_1
Xhold189 _0321_ VPWR VGND net231 sg13g2_dlygate4sd3_1
Xfanout603 _1119_ net603 VPWR VGND sg13g2_buf_8
Xfanout614 _1137_ net614 VPWR VGND sg13g2_buf_8
Xhold178 _0072_ VPWR VGND net220 sg13g2_dlygate4sd3_1
X_4377_ net730 VGND VPWR _0379_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[7\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
Xfanout636 _1061_ net636 VPWR VGND sg13g2_buf_8
X_3328_ net423 net569 _1379_ VPWR VGND sg13g2_nor2_1
Xfanout647 net658 net647 VPWR VGND sg13g2_buf_8
Xfanout658 net701 net658 VPWR VGND sg13g2_buf_8
Xfanout625 _1488_ net625 VPWR VGND sg13g2_buf_2
Xfanout669 net671 net669 VPWR VGND sg13g2_buf_8
X_3259_ net818 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[21\]
+ _1326_ VPWR VGND sg13g2_nor2_1
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_22_461 VPWR VGND sg13g2_fill_1
XFILLER_10_612 VPWR VGND sg13g2_fill_2
XFILLER_2_844 VPWR VGND sg13g2_decap_8
Xhold690 _0384_ VPWR VGND net1008 sg13g2_dlygate4sd3_1
XFILLER_1_365 VPWR VGND sg13g2_decap_8
XFILLER_45_531 VPWR VGND sg13g2_fill_2
XFILLER_17_277 VPWR VGND sg13g2_fill_2
XFILLER_14_995 VPWR VGND sg13g2_decap_8
XFILLER_9_454 VPWR VGND sg13g2_decap_4
X_2630_ net847 net413 _0905_ VPWR VGND sg13g2_nor2_2
XFILLER_9_498 VPWR VGND sg13g2_decap_4
X_2561_ _0850_ net779 _0705_ VPWR VGND sg13g2_nand2_1
X_2492_ _0480_ _0788_ _0789_ VPWR VGND sg13g2_nor2_1
X_4300_ net668 VGND VPWR _0302_ u_usb_cdc.bulk_out_nak[0] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4231_ net639 VGND VPWR net194 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[67\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
X_4162_ net673 VGND VPWR net281 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[2\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_2
X_4093_ net655 VGND VPWR net254 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[13\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3113_ VGND VPWR _1168_ net604 _0215_ _1212_ sg13g2_a21oi_1
X_3044_ _1173_ net755 net630 VPWR VGND sg13g2_nand2_1
XFILLER_23_203 VPWR VGND sg13g2_fill_1
XFILLER_36_564 VPWR VGND sg13g2_decap_8
X_3946_ _1835_ _1836_ _1834_ _1837_ VPWR VGND sg13g2_nand3_1
XFILLER_17_1001 VPWR VGND sg13g2_decap_8
X_3877_ VGND VPWR u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] _1788_ _1792_ net294
+ sg13g2_a21oi_1
XFILLER_20_976 VPWR VGND sg13g2_fill_2
X_2828_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net442 _1058_ _0084_ VPWR VGND sg13g2_mux2_1
X_2759_ net745 VPWR _1005_ VGND net832 _1004_ sg13g2_o21ai_1
X_4429_ net732 VGND VPWR net12 u_usb_cdc.u_sie.u_phy_rx.dn_q\[2\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_47_807 VPWR VGND sg13g2_decap_8
XFILLER_27_531 VPWR VGND sg13g2_fill_1
XFILLER_14_236 VPWR VGND sg13g2_fill_1
XFILLER_42_589 VPWR VGND sg13g2_fill_2
XFILLER_10_486 VPWR VGND sg13g2_fill_1
XFILLER_11_987 VPWR VGND sg13g2_decap_8
XFILLER_13_61 VPWR VGND sg13g2_fill_1
XFILLER_7_969 VPWR VGND sg13g2_decap_8
XFILLER_2_641 VPWR VGND sg13g2_decap_8
XFILLER_46_851 VPWR VGND sg13g2_decap_8
XFILLER_33_545 VPWR VGND sg13g2_decap_8
XFILLER_21_707 VPWR VGND sg13g2_fill_2
X_3800_ _0450_ VPWR _1735_ VGND u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] net515 sg13g2_o21ai_1
X_3731_ _1691_ VPWR _0354_ VGND _1900_ net598 sg13g2_o21ai_1
X_3662_ _1630_ _1632_ net789 _1633_ VPWR VGND sg13g2_nand3_1
X_3593_ _1566_ VPWR _1567_ VGND net789 _1561_ sg13g2_o21ai_1
X_2613_ net764 _0873_ _0890_ _0893_ VPWR VGND sg13g2_nor3_1
X_2544_ _0718_ _0835_ _0715_ _0836_ VPWR VGND sg13g2_nand3_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2475_ _0772_ _0662_ _0771_ VPWR VGND sg13g2_nand2_1
X_4214_ net647 VGND VPWR net277 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[50\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_4145_ net653 VGND VPWR net431 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[65\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4076_ net648 VGND VPWR _0079_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3027_ _1160_ VPWR _0180_ VGND net821 _1161_ sg13g2_o21ai_1
XFILLER_24_545 VPWR VGND sg13g2_decap_8
XFILLER_34_49 VPWR VGND sg13g2_fill_2
XFILLER_24_589 VPWR VGND sg13g2_fill_1
X_3929_ _1820_ _1821_ _1991_ _1822_ VPWR VGND sg13g2_nand3_1
XFILLER_4_928 VPWR VGND sg13g2_decap_8
XFILLER_3_427 VPWR VGND sg13g2_fill_1
XFILLER_3_416 VPWR VGND sg13g2_decap_8
XFILLER_27_383 VPWR VGND sg13g2_decap_4
XFILLER_43_887 VPWR VGND sg13g2_decap_8
XFILLER_30_526 VPWR VGND sg13g2_fill_2
XFILLER_7_733 VPWR VGND sg13g2_decap_8
XFILLER_6_265 VPWR VGND sg13g2_fill_1
XFILLER_40_92 VPWR VGND sg13g2_decap_4
XFILLER_3_983 VPWR VGND sg13g2_decap_8
X_2260_ VGND VPWR _0562_ net841 net767 sg13g2_or2_1
X_2191_ _0489_ _0490_ _0492_ _0493_ VPWR VGND sg13g2_mux2_1
XFILLER_37_103 VPWR VGND sg13g2_decap_4
XFILLER_38_637 VPWR VGND sg13g2_decap_8
XFILLER_19_851 VPWR VGND sg13g2_fill_2
XFILLER_37_125 VPWR VGND sg13g2_fill_2
XFILLER_19_884 VPWR VGND sg13g2_decap_8
XFILLER_33_320 VPWR VGND sg13g2_decap_8
XFILLER_21_526 VPWR VGND sg13g2_fill_2
X_3714_ _1665_ VPWR _0346_ VGND _1681_ _1682_ sg13g2_o21ai_1
X_3645_ _1616_ net771 _1617_ VPWR VGND sg13g2_nor2b_1
X_3576_ VGND VPWR _1549_ _1550_ _1551_ _1503_ sg13g2_a21oi_1
X_2527_ u_usb_cdc.u_ctrl_endp.rec_q\[1\] _0698_ _1926_ _0822_ VPWR VGND net618 sg13g2_nand4_1
X_2458_ u_usb_cdc.u_ctrl_endp.req_q\[1\] u_usb_cdc.u_ctrl_endp.req_q\[9\] _0747_ _0755_
+ VPWR VGND sg13g2_nor3_1
XFILLER_29_16 VPWR VGND sg13g2_decap_8
Xhold38 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[47\] VPWR VGND
+ net80 sg13g2_dlygate4sd3_1
Xhold16 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[27\] VPWR VGND
+ net58 sg13g2_dlygate4sd3_1
Xhold27 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[12\] VPWR VGND
+ net69 sg13g2_dlygate4sd3_1
Xhold49 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[15\] VPWR VGND
+ net91 sg13g2_dlygate4sd3_1
X_2389_ VPWR _0689_ _0688_ VGND sg13g2_inv_1
XFILLER_21_1019 VPWR VGND sg13g2_decap_4
X_4128_ net649 VGND VPWR net156 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[48\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_16_309 VPWR VGND sg13g2_fill_1
X_4059_ net731 VGND VPWR _0031_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[3\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
XFILLER_37_670 VPWR VGND sg13g2_decap_8
XFILLER_24_320 VPWR VGND sg13g2_decap_8
XFILLER_37_681 VPWR VGND sg13g2_fill_2
XFILLER_24_342 VPWR VGND sg13g2_decap_4
XFILLER_25_876 VPWR VGND sg13g2_decap_8
XFILLER_25_887 VPWR VGND sg13g2_fill_1
XFILLER_24_364 VPWR VGND sg13g2_fill_1
XFILLER_40_879 VPWR VGND sg13g2_decap_8
XFILLER_40_868 VPWR VGND sg13g2_fill_2
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_0_920 VPWR VGND sg13g2_decap_8
XFILLER_48_924 VPWR VGND sg13g2_decap_8
XFILLER_0_997 VPWR VGND sg13g2_decap_8
XFILLER_19_169 VPWR VGND sg13g2_fill_1
XFILLER_15_375 VPWR VGND sg13g2_decap_8
XFILLER_31_846 VPWR VGND sg13g2_decap_4
XFILLER_7_530 VPWR VGND sg13g2_fill_1
XFILLER_7_552 VPWR VGND sg13g2_decap_8
Xhold508 u_usb_cdc.u_ctrl_endp.state_q\[1\] VPWR VGND net550 sg13g2_dlygate4sd3_1
X_3430_ _1444_ net951 _1441_ VPWR VGND sg13g2_xnor2_1
Xhold519 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] VPWR VGND net561 sg13g2_dlygate4sd3_1
X_3361_ net364 net571 _1395_ VPWR VGND sg13g2_nor2_1
XFILLER_3_780 VPWR VGND sg13g2_decap_8
X_2312_ _1910_ _0563_ _0570_ _0612_ _0613_ VPWR VGND sg13g2_nor4_1
X_3292_ net960 _1271_ _1352_ _0254_ VPWR VGND sg13g2_mux2_1
X_2243_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] u_usb_cdc.u_ctrl_endp.req_q\[2\] _0545_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_39_924 VPWR VGND sg13g2_decap_8
X_2174_ _0476_ _0472_ _0475_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_445 VPWR VGND sg13g2_fill_2
XFILLER_38_478 VPWR VGND sg13g2_fill_1
X_3628_ _1592_ VPWR _1601_ VGND _1597_ _1600_ sg13g2_o21ai_1
Xoutput39 net39 usb_dp_en_o VPWR VGND sg13g2_buf_1
Xoutput28 net28 uio_out[6] VPWR VGND sg13g2_buf_1
Xoutput17 net17 uio_oe[3] VPWR VGND sg13g2_buf_1
X_3559_ VGND VPWR net799 _1968_ _1534_ net792 sg13g2_a21oi_1
XFILLER_0_249 VPWR VGND sg13g2_decap_8
XFILLER_5_1002 VPWR VGND sg13g2_decap_8
XFILLER_29_401 VPWR VGND sg13g2_decap_4
XFILLER_45_905 VPWR VGND sg13g2_decap_8
XFILLER_17_618 VPWR VGND sg13g2_decap_8
XFILLER_29_478 VPWR VGND sg13g2_fill_2
XFILLER_40_632 VPWR VGND sg13g2_decap_8
XFILLER_8_305 VPWR VGND sg13g2_fill_2
XFILLER_48_721 VPWR VGND sg13g2_decap_8
XFILLER_0_794 VPWR VGND sg13g2_decap_8
XFILLER_48_798 VPWR VGND sg13g2_decap_8
XFILLER_35_426 VPWR VGND sg13g2_decap_8
XFILLER_35_448 VPWR VGND sg13g2_fill_1
X_2930_ _1112_ VPWR _0132_ VGND net707 _1085_ sg13g2_o21ai_1
X_2861_ _1078_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ net636 VPWR VGND sg13g2_nand2_1
XFILLER_7_30 VPWR VGND sg13g2_decap_4
X_2792_ _1034_ net702 VPWR VGND net829 sg13g2_nand2b_2
XFILLER_8_861 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_fill_1
Xhold305 _1461_ VPWR VGND net347 sg13g2_dlygate4sd3_1
Xhold316 _1796_ VPWR VGND net358 sg13g2_dlygate4sd3_1
Xhold338 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[6\] VPWR VGND
+ net380 sg13g2_dlygate4sd3_1
Xhold349 u_usb_cdc.u_ctrl_endp.addr_dd\[1\] VPWR VGND net391 sg13g2_dlygate4sd3_1
X_3413_ _1431_ net783 _1424_ VPWR VGND sg13g2_nand2_1
Xhold327 _0428_ VPWR VGND net369 sg13g2_dlygate4sd3_1
Xfanout807 net808 net807 VPWR VGND sg13g2_buf_8
X_4393_ net726 VGND VPWR net298 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[14\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_3344_ net865 net458 _1384_ _0273_ VPWR VGND sg13g2_mux2_1
Xfanout818 net819 net818 VPWR VGND sg13g2_buf_8
Xfanout829 net561 net829 VPWR VGND sg13g2_buf_8
X_3275_ VPWR VGND _1336_ net807 _1340_ net810 _1341_ _1339_ sg13g2_a221oi_1
X_2226_ _0500_ _0514_ _0516_ _0527_ _0528_ VPWR VGND sg13g2_and4_1
XFILLER_39_787 VPWR VGND sg13g2_fill_1
X_2157_ _0459_ net752 u_usb_cdc.addr\[6\] VPWR VGND sg13g2_xnor2_1
XFILLER_26_39 VPWR VGND sg13g2_decap_4
X_2088_ _1966_ net310 VPWR VGND sg13g2_inv_2
XFILLER_35_971 VPWR VGND sg13g2_decap_8
XFILLER_34_492 VPWR VGND sg13g2_fill_1
XFILLER_22_654 VPWR VGND sg13g2_fill_2
XFILLER_1_547 VPWR VGND sg13g2_decap_8
XFILLER_45_757 VPWR VGND sg13g2_fill_2
XFILLER_16_83 VPWR VGND sg13g2_fill_2
XFILLER_41_996 VPWR VGND sg13g2_decap_8
XFILLER_9_658 VPWR VGND sg13g2_decap_8
XFILLER_12_175 VPWR VGND sg13g2_fill_2
XFILLER_8_179 VPWR VGND sg13g2_fill_1
XFILLER_5_820 VPWR VGND sg13g2_decap_8
XFILLER_5_897 VPWR VGND sg13g2_decap_8
XFILLER_0_591 VPWR VGND sg13g2_decap_8
X_3060_ net708 _1149_ net735 _1184_ VPWR VGND _1183_ sg13g2_nand4_1
XFILLER_48_551 VPWR VGND sg13g2_decap_8
XFILLER_35_201 VPWR VGND sg13g2_fill_2
XFILLER_36_724 VPWR VGND sg13g2_decap_8
XFILLER_36_735 VPWR VGND sg13g2_fill_1
XFILLER_35_223 VPWR VGND sg13g2_decap_4
X_3962_ _1851_ net274 net621 VPWR VGND sg13g2_nand2_1
X_3893_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] net973 net704 _0407_ VPWR VGND sg13g2_mux2_1
XFILLER_32_985 VPWR VGND sg13g2_decap_8
X_2913_ _1103_ VPWR _0124_ VGND _1066_ net615 sg13g2_o21ai_1
X_2844_ _1065_ VPWR _0092_ VGND net616 _1066_ sg13g2_o21ai_1
X_2775_ _1013_ _1018_ _1019_ _1020_ VPWR VGND sg13g2_nor3_1
Xhold135 _0195_ VPWR VGND net177 sg13g2_dlygate4sd3_1
Xhold102 _0238_ VPWR VGND net144 sg13g2_dlygate4sd3_1
Xhold113 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[48\] VPWR VGND
+ net155 sg13g2_dlygate4sd3_1
Xhold124 _0437_ VPWR VGND net166 sg13g2_dlygate4sd3_1
Xhold168 _0058_ VPWR VGND net210 sg13g2_dlygate4sd3_1
Xhold157 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[57\] VPWR
+ VGND net199 sg13g2_dlygate4sd3_1
Xhold146 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[33\] VPWR
+ VGND net188 sg13g2_dlygate4sd3_1
X_4445_ net726 VGND VPWR _0041_ u_usb_cdc.clk_gate_q clknet_leaf_40_clk sg13g2_dfrbpq_2
Xfanout615 _1099_ net615 VPWR VGND sg13g2_buf_8
Xfanout604 net605 net604 VPWR VGND sg13g2_buf_8
Xhold179 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[15\] VPWR
+ VGND net221 sg13g2_dlygate4sd3_1
X_4376_ net730 VGND VPWR _0378_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[6\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
X_3327_ VGND VPWR _1894_ net569 _0263_ _1378_ sg13g2_a21oi_1
Xfanout648 net649 net648 VPWR VGND sg13g2_buf_8
Xfanout637 net638 net637 VPWR VGND sg13g2_buf_8
Xfanout626 _1360_ net626 VPWR VGND sg13g2_buf_8
Xfanout659 net661 net659 VPWR VGND sg13g2_buf_8
XFILLER_2_1005 VPWR VGND sg13g2_decap_8
X_3258_ net818 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[37\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[45\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[53\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[61\] net811 _1325_
+ VPWR VGND sg13g2_mux4_1
XFILLER_37_27 VPWR VGND sg13g2_decap_4
X_2209_ _0511_ u_usb_cdc.u_sie.crc16_q\[14\] net764 VPWR VGND sg13g2_xnor2_1
X_3189_ net578 net1015 _1263_ _0240_ VPWR VGND sg13g2_a21o_1
XFILLER_14_418 VPWR VGND sg13g2_fill_1
XFILLER_26_267 VPWR VGND sg13g2_decap_8
XFILLER_35_790 VPWR VGND sg13g2_fill_1
XFILLER_5_116 VPWR VGND sg13g2_fill_2
XFILLER_5_138 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
Xhold680 _0159_ VPWR VGND net998 sg13g2_dlygate4sd3_1
Xhold691 u_usb_cdc.u_sie.pid_q\[2\] VPWR VGND net1009 sg13g2_dlygate4sd3_1
XFILLER_18_702 VPWR VGND sg13g2_decap_4
XFILLER_18_724 VPWR VGND sg13g2_fill_2
XFILLER_27_93 VPWR VGND sg13g2_fill_1
XFILLER_14_974 VPWR VGND sg13g2_decap_4
X_2560_ u_usb_cdc.u_ctrl_endp.max_length_q\[6\] _0847_ _0848_ _0849_ VPWR VGND sg13g2_nor3_1
X_2491_ u_usb_cdc.sie_out_data\[2\] _0707_ net719 _0788_ VPWR VGND sg13g2_nand3_1
XFILLER_5_694 VPWR VGND sg13g2_decap_8
X_4230_ net639 VGND VPWR net121 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[66\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4161_ net672 VGND VPWR net928 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[1\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_2
X_3112_ net362 net604 _1212_ VPWR VGND sg13g2_nor2_1
X_4092_ net669 VGND VPWR net70 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[12\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_49_893 VPWR VGND sg13g2_decap_8
X_3043_ VGND VPWR net611 _1172_ _0185_ _1171_ sg13g2_a21oi_1
XFILLER_36_521 VPWR VGND sg13g2_fill_2
X_3945_ _1836_ u_usb_cdc.u_sie.data_q\[3\] net834 u_usb_cdc.u_sie.pid_q\[3\] net830
+ VPWR VGND sg13g2_a22oi_1
X_3876_ VGND VPWR _1788_ _1790_ _1791_ net704 sg13g2_a21oi_1
X_2827_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net378 _1058_ _0083_ VPWR VGND sg13g2_mux2_1
X_2758_ net766 _1003_ _1004_ VPWR VGND sg13g2_nor2_1
X_2689_ VGND VPWR _1961_ _0949_ _0035_ _0952_ sg13g2_a21oi_1
X_4428_ net732 VGND VPWR net43 u_usb_cdc.u_sie.u_phy_rx.dn_q\[1\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_48_37 VPWR VGND sg13g2_fill_1
XFILLER_24_1017 VPWR VGND sg13g2_decap_8
X_4359_ net648 VGND VPWR net504 net20 clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_42_513 VPWR VGND sg13g2_fill_2
XFILLER_11_966 VPWR VGND sg13g2_decap_8
XFILLER_10_476 VPWR VGND sg13g2_fill_2
XFILLER_7_948 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_fill_1
XFILLER_2_620 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_8
XFILLER_37_307 VPWR VGND sg13g2_decap_8
XFILLER_46_830 VPWR VGND sg13g2_decap_8
X_3730_ net590 _1683_ net919 _1691_ VPWR VGND sg13g2_nand3_1
X_3661_ _1632_ net791 _1631_ VPWR VGND sg13g2_nand2_1
X_3592_ _1566_ _1563_ _1565_ VPWR VGND sg13g2_nand2_1
X_2612_ _0871_ VPWR _0021_ VGND _0873_ _0892_ sg13g2_o21ai_1
X_2543_ net574 VPWR _0835_ VGND _0674_ _0675_ sg13g2_o21ai_1
XFILLER_47_1017 VPWR VGND sg13g2_decap_8
X_2474_ _0770_ VPWR _0771_ VGND _1931_ _0767_ sg13g2_o21ai_1
X_4213_ net659 VGND VPWR net417 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[49\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_29_819 VPWR VGND sg13g2_fill_1
X_4144_ net653 VGND VPWR net451 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[64\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_28_318 VPWR VGND sg13g2_decap_4
XFILLER_49_690 VPWR VGND sg13g2_decap_8
X_4075_ net648 VGND VPWR _0078_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3026_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[0\] _1150_
+ net753 _1161_ VPWR VGND sg13g2_nand3_1
XFILLER_24_502 VPWR VGND sg13g2_decap_8
XFILLER_24_568 VPWR VGND sg13g2_fill_2
X_3928_ _1821_ _1953_ net831 net765 net834 VPWR VGND sg13g2_a22oi_1
X_3859_ net297 _1776_ _1779_ VPWR VGND sg13g2_and2_1
XFILLER_4_907 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_8_1022 VPWR VGND sg13g2_decap_8
XFILLER_27_373 VPWR VGND sg13g2_decap_4
XFILLER_43_866 VPWR VGND sg13g2_decap_8
XFILLER_7_712 VPWR VGND sg13g2_decap_8
XFILLER_7_789 VPWR VGND sg13g2_decap_8
XFILLER_3_962 VPWR VGND sg13g2_decap_8
XFILLER_2_483 VPWR VGND sg13g2_decap_8
X_2190_ _0476_ u_usb_cdc.u_sie.data_q\[5\] _0492_ VPWR VGND sg13g2_xor2_1
XFILLER_1_21 VPWR VGND sg13g2_fill_2
XFILLER_19_841 VPWR VGND sg13g2_fill_2
XFILLER_46_682 VPWR VGND sg13g2_decap_8
XFILLER_34_877 VPWR VGND sg13g2_fill_2
XFILLER_33_387 VPWR VGND sg13g2_decap_4
XFILLER_34_899 VPWR VGND sg13g2_decap_4
XFILLER_14_1016 VPWR VGND sg13g2_decap_8
XFILLER_14_1027 VPWR VGND sg13g2_fill_2
X_3713_ net597 VPWR _1682_ VGND net999 net624 sg13g2_o21ai_1
X_3644_ net781 _0549_ _0670_ _1616_ VPWR VGND sg13g2_nor3_1
X_3575_ _0542_ _0664_ _1550_ VPWR VGND net776 sg13g2_nand3b_1
XFILLER_0_409 VPWR VGND sg13g2_decap_8
X_2526_ _0679_ _0680_ _0821_ VPWR VGND sg13g2_nor2_1
X_2457_ _0754_ _0752_ _0753_ VPWR VGND sg13g2_nand2_1
XFILLER_29_39 VPWR VGND sg13g2_fill_2
Xhold28 _0095_ VPWR VGND net70 sg13g2_dlygate4sd3_1
Xhold17 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[55\] VPWR VGND
+ net59 sg13g2_dlygate4sd3_1
Xhold39 _0130_ VPWR VGND net81 sg13g2_dlygate4sd3_1
X_2388_ _0542_ _0654_ _0688_ VPWR VGND sg13g2_nor2_2
XFILLER_29_616 VPWR VGND sg13g2_fill_2
XFILLER_29_638 VPWR VGND sg13g2_fill_2
X_4127_ net669 VGND VPWR net81 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[47\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_4058_ net731 VGND VPWR net1013 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
XFILLER_45_49 VPWR VGND sg13g2_fill_1
X_3009_ _1149_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\]
+ _1148_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_704 VPWR VGND sg13g2_decap_8
XFILLER_3_203 VPWR VGND sg13g2_fill_2
XFILLER_48_903 VPWR VGND sg13g2_decap_8
XFILLER_0_976 VPWR VGND sg13g2_decap_8
XFILLER_16_833 VPWR VGND sg13g2_fill_2
XFILLER_34_107 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_54_clk clknet_3_0__leaf_clk clknet_leaf_54_clk VPWR VGND sg13g2_buf_8
XFILLER_43_696 VPWR VGND sg13g2_fill_2
XFILLER_30_313 VPWR VGND sg13g2_decap_8
Xhold509 _0011_ VPWR VGND net551 sg13g2_dlygate4sd3_1
X_3360_ VGND VPWR _1898_ net571 _0280_ _1394_ sg13g2_a21oi_1
X_2311_ u_usb_cdc.u_sie.in_byte_q\[3\] _1989_ _0611_ _0612_ VPWR VGND sg13g2_nor3_1
X_3291_ net983 _1265_ _1352_ _0253_ VPWR VGND sg13g2_mux2_1
XFILLER_32_4 VPWR VGND sg13g2_decap_4
XFILLER_39_903 VPWR VGND sg13g2_decap_8
X_2242_ net770 net773 _0544_ VPWR VGND sg13g2_nor2b_2
XFILLER_38_413 VPWR VGND sg13g2_fill_1
X_2173_ _0475_ _0473_ _0474_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_424 VPWR VGND sg13g2_fill_2
XFILLER_25_118 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_45_clk clknet_3_4__leaf_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
XFILLER_18_192 VPWR VGND sg13g2_fill_1
XFILLER_33_140 VPWR VGND sg13g2_fill_2
XFILLER_21_324 VPWR VGND sg13g2_fill_1
X_3627_ _1599_ VPWR _1600_ VGND net771 _1544_ sg13g2_o21ai_1
Xoutput29 net29 uo_out[0] VPWR VGND sg13g2_buf_1
Xoutput18 net18 uio_oe[4] VPWR VGND sg13g2_buf_1
X_3558_ net797 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[1\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[9\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[17\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[25\]
+ net792 _1533_ VPWR VGND sg13g2_mux4_1
X_2509_ VGND VPWR _0801_ _0802_ _0806_ _0798_ sg13g2_a21oi_1
XFILLER_1_729 VPWR VGND sg13g2_decap_8
X_3489_ net835 net839 _1481_ VPWR VGND sg13g2_nor2_1
XFILLER_29_424 VPWR VGND sg13g2_fill_1
XFILLER_38_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_36_clk clknet_3_4__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_37_490 VPWR VGND sg13g2_fill_2
XFILLER_25_685 VPWR VGND sg13g2_decap_4
XFILLER_40_611 VPWR VGND sg13g2_fill_1
XFILLER_12_324 VPWR VGND sg13g2_fill_1
XFILLER_13_836 VPWR VGND sg13g2_fill_1
XFILLER_40_655 VPWR VGND sg13g2_fill_2
XFILLER_9_829 VPWR VGND sg13g2_fill_1
XFILLER_40_699 VPWR VGND sg13g2_decap_8
XFILLER_8_339 VPWR VGND sg13g2_decap_8
XFILLER_43_1020 VPWR VGND sg13g2_decap_8
XFILLER_0_773 VPWR VGND sg13g2_decap_8
XFILLER_47_221 VPWR VGND sg13g2_decap_8
XFILLER_48_777 VPWR VGND sg13g2_decap_8
XFILLER_47_232 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_27_clk clknet_3_6__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_44_983 VPWR VGND sg13g2_decap_8
XFILLER_43_482 VPWR VGND sg13g2_decap_4
X_2860_ _1077_ net91 _1059_ VPWR VGND sg13g2_nand2_1
XFILLER_31_655 VPWR VGND sg13g2_decap_4
X_2791_ net829 _1993_ _1033_ VPWR VGND sg13g2_nor2_1
XFILLER_11_1008 VPWR VGND sg13g2_decap_8
XFILLER_7_372 VPWR VGND sg13g2_fill_2
XFILLER_7_86 VPWR VGND sg13g2_fill_1
Xhold306 _0314_ VPWR VGND net348 sg13g2_dlygate4sd3_1
Xhold317 _0403_ VPWR VGND net359 sg13g2_dlygate4sd3_1
Xhold339 _0089_ VPWR VGND net381 sg13g2_dlygate4sd3_1
Xhold328 net19 VPWR VGND net370 sg13g2_dlygate4sd3_1
X_3412_ _1428_ VPWR _0296_ VGND _1426_ _1430_ sg13g2_o21ai_1
X_4392_ net726 VGND VPWR net367 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[13\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_3343_ net896 net384 _1384_ _0272_ VPWR VGND sg13g2_mux2_1
Xfanout819 net1054 net819 VPWR VGND sg13g2_buf_8
Xfanout808 net1024 net808 VPWR VGND sg13g2_buf_8
X_3274_ VGND VPWR net813 _1979_ _1340_ net809 sg13g2_a21oi_1
X_2225_ _0519_ _0520_ _0522_ _0526_ _0527_ VPWR VGND sg13g2_nor4_1
XFILLER_38_221 VPWR VGND sg13g2_fill_2
X_2156_ _0458_ net753 u_usb_cdc.addr\[5\] VPWR VGND sg13g2_xnor2_1
X_2087_ VPWR _0039_ net48 VGND sg13g2_inv_1
XFILLER_35_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_3_3__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_21_143 VPWR VGND sg13g2_fill_1
X_2989_ _1137_ _1136_ VPWR VGND net630 sg13g2_nand2b_2
XFILLER_22_699 VPWR VGND sg13g2_decap_8
XFILLER_5_309 VPWR VGND sg13g2_fill_2
XFILLER_1_526 VPWR VGND sg13g2_decap_8
XFILLER_49_519 VPWR VGND sg13g2_decap_8
XFILLER_45_736 VPWR VGND sg13g2_decap_8
XFILLER_29_265 VPWR VGND sg13g2_decap_8
XFILLER_45_769 VPWR VGND sg13g2_decap_8
XFILLER_16_40 VPWR VGND sg13g2_fill_2
XFILLER_26_994 VPWR VGND sg13g2_decap_8
XFILLER_13_611 VPWR VGND sg13g2_decap_8
XFILLER_25_482 VPWR VGND sg13g2_fill_1
XFILLER_41_975 VPWR VGND sg13g2_decap_8
XFILLER_34_1008 VPWR VGND sg13g2_decap_8
XFILLER_40_430 VPWR VGND sg13g2_decap_4
XFILLER_40_441 VPWR VGND sg13g2_fill_1
XFILLER_9_648 VPWR VGND sg13g2_fill_1
XFILLER_40_474 VPWR VGND sg13g2_decap_4
XFILLER_5_876 VPWR VGND sg13g2_decap_8
XFILLER_0_570 VPWR VGND sg13g2_decap_8
XFILLER_48_530 VPWR VGND sg13g2_decap_8
XFILLER_36_703 VPWR VGND sg13g2_decap_4
X_3961_ _0425_ _1849_ _1850_ net621 _1977_ VPWR VGND sg13g2_a22oi_1
XFILLER_17_972 VPWR VGND sg13g2_fill_2
XFILLER_44_791 VPWR VGND sg13g2_decap_8
XFILLER_44_780 VPWR VGND sg13g2_fill_2
X_2912_ _1103_ net73 _1101_ VPWR VGND sg13g2_nand2_1
X_3892_ VGND VPWR net744 _0973_ _0406_ net977 sg13g2_a21oi_1
XFILLER_32_964 VPWR VGND sg13g2_decap_8
XFILLER_31_485 VPWR VGND sg13g2_fill_2
X_2843_ _1066_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2774_ VGND VPWR _1907_ _1987_ _1019_ _1908_ sg13g2_a21oi_1
XFILLER_8_681 VPWR VGND sg13g2_decap_8
Xhold103 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[65\] VPWR
+ VGND net145 sg13g2_dlygate4sd3_1
Xhold125 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[61\] VPWR
+ VGND net167 sg13g2_dlygate4sd3_1
Xhold114 _0131_ VPWR VGND net156 sg13g2_dlygate4sd3_1
Xhold136 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[18\] VPWR VGND
+ net178 sg13g2_dlygate4sd3_1
Xhold158 u_usb_cdc.u_sie.addr_q\[3\] VPWR VGND net200 sg13g2_dlygate4sd3_1
Xhold147 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[17\] VPWR VGND net189 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_4__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
X_4444_ net699 VGND VPWR net334 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[2\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
Xhold169 u_usb_cdc.u_sie.u_phy_tx.data_q\[2\] VPWR VGND net211 sg13g2_dlygate4sd3_1
Xfanout605 _1211_ net605 VPWR VGND sg13g2_buf_8
X_4375_ net730 VGND VPWR _0377_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[5\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
Xfanout616 _1064_ net616 VPWR VGND sg13g2_buf_8
Xfanout627 net629 net627 VPWR VGND sg13g2_buf_8
X_3326_ net518 net569 _1378_ VPWR VGND sg13g2_nor2_1
Xfanout649 net652 net649 VPWR VGND sg13g2_buf_8
Xfanout638 _1038_ net638 VPWR VGND sg13g2_buf_8
X_3257_ _0247_ _1324_ _1323_ VPWR VGND sg13g2_nand2b_1
X_2208_ net766 net915 _0510_ VPWR VGND sg13g2_xor2_1
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
X_3188_ VGND VPWR _1261_ _1262_ _1263_ net578 sg13g2_a21oi_1
X_2139_ _1934_ _1935_ _0442_ VPWR VGND sg13g2_nor2_1
XFILLER_23_931 VPWR VGND sg13g2_fill_1
XFILLER_22_430 VPWR VGND sg13g2_decap_8
XFILLER_10_614 VPWR VGND sg13g2_fill_1
XFILLER_6_629 VPWR VGND sg13g2_decap_8
XFILLER_2_802 VPWR VGND sg13g2_decap_8
Xhold670 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] VPWR VGND net988 sg13g2_dlygate4sd3_1
Xhold681 u_usb_cdc.u_sie.rx_data\[7\] VPWR VGND net999 sg13g2_dlygate4sd3_1
XFILLER_2_879 VPWR VGND sg13g2_decap_8
Xhold692 _0368_ VPWR VGND net1010 sg13g2_dlygate4sd3_1
XFILLER_40_1012 VPWR VGND sg13g2_decap_8
XFILLER_17_202 VPWR VGND sg13g2_fill_2
XFILLER_45_555 VPWR VGND sg13g2_decap_8
XFILLER_13_441 VPWR VGND sg13g2_decap_8
XFILLER_13_452 VPWR VGND sg13g2_fill_1
XFILLER_9_478 VPWR VGND sg13g2_decap_8
XFILLER_4_150 VPWR VGND sg13g2_fill_1
X_2490_ _0777_ _0779_ _0774_ _0787_ VPWR VGND _0786_ sg13g2_nand4_1
X_4160_ net673 VGND VPWR net302 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[0\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_1_890 VPWR VGND sg13g2_decap_8
X_3111_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\] net820
+ _1964_ _1136_ _1211_ VPWR VGND sg13g2_and4_1
X_4091_ net655 VGND VPWR net138 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[11\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_49_872 VPWR VGND sg13g2_decap_8
X_3042_ _1172_ net756 net630 VPWR VGND sg13g2_nand2_2
XFILLER_36_544 VPWR VGND sg13g2_fill_2
X_3944_ _1835_ _1951_ net831 _1941_ net838 VPWR VGND sg13g2_a22oi_1
X_3875_ _1790_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] net294 VPWR VGND sg13g2_nand2_1
X_2826_ _1058_ _1040_ _1057_ VPWR VGND sg13g2_nand2_2
XFILLER_20_978 VPWR VGND sg13g2_fill_1
X_2757_ _1003_ net765 _0889_ VPWR VGND sg13g2_nand2_1
XFILLER_2_109 VPWR VGND sg13g2_fill_1
X_2688_ net342 net987 _0952_ VPWR VGND sg13g2_nor2_2
X_4427_ net731 VGND VPWR net46 u_usb_cdc.u_sie.u_phy_rx.dn_q\[0\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
X_4358_ net648 VGND VPWR net371 net19 clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4289_ net662 VGND VPWR net917 u_usb_cdc.u_ctrl_endp.max_length_q\[3\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_3309_ _1364_ net803 net795 VPWR VGND sg13g2_xnor2_1
XFILLER_11_945 VPWR VGND sg13g2_decap_8
XFILLER_22_282 VPWR VGND sg13g2_fill_2
XFILLER_22_293 VPWR VGND sg13g2_fill_1
XFILLER_7_927 VPWR VGND sg13g2_decap_8
XFILLER_6_404 VPWR VGND sg13g2_fill_2
XFILLER_2_676 VPWR VGND sg13g2_decap_8
XFILLER_46_886 VPWR VGND sg13g2_decap_8
XFILLER_18_599 VPWR VGND sg13g2_fill_2
XFILLER_14_794 VPWR VGND sg13g2_fill_1
X_3660_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[53\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[61\]
+ net797 _1631_ VPWR VGND sg13g2_mux2_1
X_3591_ VGND VPWR net791 _1564_ _1565_ _1913_ sg13g2_a21oi_1
X_2611_ _0892_ net764 _0891_ VPWR VGND sg13g2_nand2_1
XFILLER_6_982 VPWR VGND sg13g2_decap_8
X_2542_ _0009_ _0833_ _0834_ VPWR VGND sg13g2_nand2_1
X_4212_ net659 VGND VPWR net363 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[48\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_2473_ _0770_ _0769_ u_usb_cdc.u_ctrl_endp.req_q\[1\] _0710_ u_usb_cdc.u_ctrl_endp.req_q\[11\]
+ VPWR VGND sg13g2_a22oi_1
X_4143_ net668 VGND VPWR net338 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[63\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_4074_ net649 VGND VPWR _0077_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_2
X_3025_ _1160_ net225 _1146_ VPWR VGND sg13g2_nand2_1
XFILLER_37_853 VPWR VGND sg13g2_fill_1
XFILLER_37_886 VPWR VGND sg13g2_fill_1
X_3927_ _1820_ _1939_ net838 u_usb_cdc.u_sie.pid_q\[1\] net830 VPWR VGND sg13g2_a22oi_1
X_3858_ _1778_ net711 net297 VPWR VGND sg13g2_nand2_1
XFILLER_20_775 VPWR VGND sg13g2_fill_1
X_2809_ _1050_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[2\] _1049_
+ VPWR VGND sg13g2_xnor2_1
X_3789_ VPWR _0377_ net863 VGND sg13g2_inv_1
XFILLER_8_1001 VPWR VGND sg13g2_decap_8
XFILLER_27_352 VPWR VGND sg13g2_decap_8
XFILLER_43_834 VPWR VGND sg13g2_decap_8
XFILLER_28_897 VPWR VGND sg13g2_decap_8
XFILLER_30_528 VPWR VGND sg13g2_fill_1
XFILLER_7_768 VPWR VGND sg13g2_decap_8
XFILLER_6_289 VPWR VGND sg13g2_fill_2
XFILLER_3_941 VPWR VGND sg13g2_decap_8
XFILLER_2_462 VPWR VGND sg13g2_decap_8
XFILLER_46_694 VPWR VGND sg13g2_decap_4
X_3712_ _1489_ _1678_ _1680_ _1681_ VPWR VGND sg13g2_nor3_1
X_3643_ _1615_ _1609_ _1614_ net626 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[68\]
+ VPWR VGND sg13g2_a22oi_1
X_3574_ net776 VPWR _1549_ VGND net781 _1429_ sg13g2_o21ai_1
X_2525_ _0814_ _0819_ _0719_ _0820_ VPWR VGND sg13g2_nand3_1
X_2456_ u_usb_cdc.u_ctrl_endp.req_q\[4\] net842 u_usb_cdc.u_ctrl_endp.req_q\[7\] _0753_
+ VPWR VGND sg13g2_nor3_1
Xhold29 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[46\] VPWR VGND
+ net71 sg13g2_dlygate4sd3_1
Xhold18 _0138_ VPWR VGND net60 sg13g2_dlygate4sd3_1
X_4126_ net670 VGND VPWR net72 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[46\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2387_ net586 net584 net619 _0686_ _0687_ VPWR VGND sg13g2_nor4_1
X_4057_ net728 VGND VPWR net893 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[1\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_3008_ net822 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\]
+ net820 _1148_ VPWR VGND sg13g2_nor3_2
XFILLER_25_834 VPWR VGND sg13g2_decap_4
XFILLER_40_826 VPWR VGND sg13g2_decap_4
XFILLER_40_848 VPWR VGND sg13g2_fill_2
XFILLER_10_31 VPWR VGND sg13g2_fill_2
XFILLER_0_955 VPWR VGND sg13g2_decap_8
XFILLER_48_959 VPWR VGND sg13g2_decap_8
XFILLER_19_116 VPWR VGND sg13g2_fill_1
XFILLER_47_469 VPWR VGND sg13g2_fill_2
XFILLER_28_650 VPWR VGND sg13g2_decap_8
XFILLER_15_322 VPWR VGND sg13g2_decap_8
XFILLER_37_1017 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_7_521 VPWR VGND sg13g2_fill_1
XFILLER_7_510 VPWR VGND sg13g2_decap_8
XFILLER_7_598 VPWR VGND sg13g2_decap_4
X_2310_ net289 net230 net319 _0611_ VPWR VGND sg13g2_nand3_1
X_3290_ net968 _1260_ _1352_ _0252_ VPWR VGND sg13g2_mux2_1
X_2241_ net786 net782 net779 _0543_ VPWR VGND sg13g2_nor3_1
X_2172_ _0474_ u_usb_cdc.sie_out_data\[0\] net762 VPWR VGND sg13g2_xnor2_1
XFILLER_39_959 VPWR VGND sg13g2_decap_8
XFILLER_33_152 VPWR VGND sg13g2_fill_1
XFILLER_34_697 VPWR VGND sg13g2_fill_1
X_3626_ _1502_ VPWR _1599_ VGND _1542_ _1598_ sg13g2_o21ai_1
XFILLER_1_708 VPWR VGND sg13g2_decap_8
Xoutput19 net19 uio_oe[5] VPWR VGND sg13g2_buf_1
X_3557_ _1532_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[65\] net626
+ VPWR VGND sg13g2_nand2_1
X_2508_ _0726_ _0802_ _0805_ VPWR VGND sg13g2_nor2_1
X_3488_ _1479_ VPWR _0322_ VGND _0894_ _1480_ sg13g2_o21ai_1
X_2439_ net884 _0734_ _0736_ _0737_ VPWR VGND sg13g2_or3_1
XFILLER_29_414 VPWR VGND sg13g2_fill_1
X_4109_ net656 VGND VPWR net411 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[29\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_38_970 VPWR VGND sg13g2_decap_8
XFILLER_37_480 VPWR VGND sg13g2_fill_1
XFILLER_24_130 VPWR VGND sg13g2_fill_1
XFILLER_25_675 VPWR VGND sg13g2_decap_4
XFILLER_8_307 VPWR VGND sg13g2_fill_1
XFILLER_0_752 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_fill_2
XFILLER_44_962 VPWR VGND sg13g2_decap_8
XFILLER_30_188 VPWR VGND sg13g2_decap_8
X_2790_ _1032_ net308 net713 VPWR VGND sg13g2_nand2_1
Xhold307 u_usb_cdc.u_sie.crc16_q\[6\] VPWR VGND net349 sg13g2_dlygate4sd3_1
XFILLER_8_896 VPWR VGND sg13g2_decap_8
X_4460_ net37 net39 VPWR VGND sg13g2_buf_1
X_4391_ net726 VGND VPWR _0393_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[12\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_3411_ _1430_ _0549_ _0661_ VPWR VGND sg13g2_nand2_1
Xhold329 _0360_ VPWR VGND net371 sg13g2_dlygate4sd3_1
Xhold318 _0056_ VPWR VGND net360 sg13g2_dlygate4sd3_1
X_3342_ net905 net510 _1384_ _0271_ VPWR VGND sg13g2_mux2_1
Xfanout809 net810 net809 VPWR VGND sg13g2_buf_8
X_3273_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[22\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[30\]
+ net813 _1339_ VPWR VGND sg13g2_mux2_1
X_2224_ _0523_ _0525_ _0507_ _0526_ VPWR VGND sg13g2_nand3_1
X_2155_ _0452_ _0454_ net352 _0457_ _0064_ VPWR VGND sg13g2_nor4_1
X_2086_ _1965_ net826 VPWR VGND sg13g2_inv_2
X_2988_ net714 net822 _1136_ VPWR VGND sg13g2_nor2_2
XFILLER_21_188 VPWR VGND sg13g2_fill_2
X_3609_ _1582_ net1011 net593 VPWR VGND sg13g2_nand2_1
XFILLER_1_505 VPWR VGND sg13g2_decap_8
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
XFILLER_45_715 VPWR VGND sg13g2_decap_8
XFILLER_45_759 VPWR VGND sg13g2_fill_1
XFILLER_26_940 VPWR VGND sg13g2_fill_1
XFILLER_16_85 VPWR VGND sg13g2_fill_1
XFILLER_41_954 VPWR VGND sg13g2_decap_8
XFILLER_9_627 VPWR VGND sg13g2_fill_1
XFILLER_5_855 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_fill_1
XFILLER_35_236 VPWR VGND sg13g2_decap_4
XFILLER_35_258 VPWR VGND sg13g2_decap_8
X_3960_ VGND VPWR net274 _1814_ _1850_ net622 sg13g2_a21oi_1
X_2911_ _1102_ VPWR _0123_ VGND _1062_ net615 sg13g2_o21ai_1
XFILLER_32_943 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
X_3891_ net746 net743 _1800_ VPWR VGND sg13g2_nor2_1
XFILLER_31_431 VPWR VGND sg13g2_decap_8
X_2842_ _1065_ net75 _1059_ VPWR VGND sg13g2_nand2_1
X_2773_ _1017_ VPWR _1018_ VGND _1966_ _0573_ sg13g2_o21ai_1
Xhold115 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[4\] VPWR VGND
+ net157 sg13g2_dlygate4sd3_1
XFILLER_7_181 VPWR VGND sg13g2_fill_1
Xhold104 _0232_ VPWR VGND net146 sg13g2_dlygate4sd3_1
Xhold126 _0228_ VPWR VGND net168 sg13g2_dlygate4sd3_1
Xhold137 _0101_ VPWR VGND net179 sg13g2_dlygate4sd3_1
Xhold159 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[31\] VPWR
+ VGND net201 sg13g2_dlygate4sd3_1
Xhold148 _0398_ VPWR VGND net190 sg13g2_dlygate4sd3_1
X_4443_ net699 VGND VPWR net317 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[1\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
Xfanout606 net607 net606 VPWR VGND sg13g2_buf_8
X_4374_ net730 VGND VPWR _0376_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[4\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
Xfanout639 net643 net639 VPWR VGND sg13g2_buf_8
Xfanout617 net618 net617 VPWR VGND sg13g2_buf_8
Xfanout628 net629 net628 VPWR VGND sg13g2_buf_1
X_3325_ _0724_ _1376_ _1377_ VPWR VGND sg13g2_nor2_2
X_3256_ _1324_ _1296_ net100 net601 net544 VPWR VGND sg13g2_a22oi_1
X_2207_ u_usb_cdc.u_sie.data_q\[4\] u_usb_cdc.u_sie.crc16_q\[11\] _0509_ VPWR VGND
+ sg13g2_xor2_1
X_3187_ _1262_ _0606_ _1260_ net968 net749 VPWR VGND sg13g2_a22oi_1
X_2138_ _0441_ _1934_ _1935_ VPWR VGND sg13g2_nand2_2
X_2069_ _1948_ net372 VPWR VGND sg13g2_inv_2
XFILLER_34_291 VPWR VGND sg13g2_decap_8
XFILLER_6_608 VPWR VGND sg13g2_decap_4
Xhold671 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[2\] VPWR VGND
+ net989 sg13g2_dlygate4sd3_1
XFILLER_2_858 VPWR VGND sg13g2_decap_8
Xhold660 _0406_ VPWR VGND net978 sg13g2_dlygate4sd3_1
Xhold682 _0060_ VPWR VGND net1000 sg13g2_dlygate4sd3_1
Xhold693 u_usb_cdc.u_sie.data_q\[3\] VPWR VGND net1011 sg13g2_dlygate4sd3_1
XFILLER_1_379 VPWR VGND sg13g2_decap_8
XFILLER_32_228 VPWR VGND sg13g2_fill_1
XFILLER_4_173 VPWR VGND sg13g2_fill_2
X_3110_ _1210_ VPWR _0214_ VGND net709 _1165_ sg13g2_o21ai_1
XFILLER_49_851 VPWR VGND sg13g2_decap_8
X_4090_ net656 VGND VPWR net192 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[10\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3041_ net321 net611 _1171_ VPWR VGND sg13g2_nor2_1
XFILLER_36_523 VPWR VGND sg13g2_fill_1
XFILLER_17_1015 VPWR VGND sg13g2_decap_8
XFILLER_23_239 VPWR VGND sg13g2_decap_4
X_3943_ _1990_ VPWR _1834_ VGND _0579_ _1018_ sg13g2_o21ai_1
X_3874_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\]
+ _1789_ VPWR VGND sg13g2_and2_1
XFILLER_31_261 VPWR VGND sg13g2_fill_1
X_2825_ net714 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] _1057_
+ VPWR VGND sg13g2_nor2_2
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_9_980 VPWR VGND sg13g2_decap_8
X_2756_ VGND VPWR net739 _0995_ _0068_ net850 sg13g2_a21oi_1
X_2687_ VPWR _0034_ net498 VGND sg13g2_inv_1
X_4426_ net725 VGND VPWR net13 u_usb_cdc.u_sie.u_phy_rx.dp_q\[2\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_4357_ net642 VGND VPWR net859 net18 clknet_leaf_3_clk sg13g2_dfrbpq_1
X_3308_ VGND VPWR _1912_ _1358_ _0259_ _1363_ sg13g2_a21oi_1
X_4288_ net666 VGND VPWR net524 u_usb_cdc.u_ctrl_endp.max_length_q\[2\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_3239_ _1307_ VPWR _1308_ VGND net812 net77 sg13g2_o21ai_1
XFILLER_27_567 VPWR VGND sg13g2_fill_2
XFILLER_11_924 VPWR VGND sg13g2_decap_8
XFILLER_22_261 VPWR VGND sg13g2_decap_8
XFILLER_7_906 VPWR VGND sg13g2_decap_8
XFILLER_6_416 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
Xhold490 _1721_ VPWR VGND net532 sg13g2_dlygate4sd3_1
XFILLER_46_865 VPWR VGND sg13g2_decap_8
XFILLER_45_353 VPWR VGND sg13g2_decap_8
XFILLER_18_567 VPWR VGND sg13g2_fill_2
XFILLER_45_364 VPWR VGND sg13g2_fill_1
XFILLER_41_570 VPWR VGND sg13g2_fill_1
X_3590_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[50\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[58\]
+ net798 _1564_ VPWR VGND sg13g2_mux2_1
X_2610_ _0882_ _0884_ _0890_ _0891_ VPWR VGND sg13g2_nor3_1
XFILLER_6_961 VPWR VGND sg13g2_decap_8
X_2541_ _0743_ _0780_ _0695_ _0834_ VPWR VGND sg13g2_nand3_1
X_2472_ VGND VPWR _1927_ _0768_ _0769_ _0767_ sg13g2_a21oi_1
X_4211_ net647 VGND VPWR net113 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[47\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
X_4142_ net672 VGND VPWR net463 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[62\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_4073_ net652 VGND VPWR _0076_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3024_ _1158_ VPWR _0179_ VGND net821 _1159_ sg13g2_o21ai_1
XFILLER_37_832 VPWR VGND sg13g2_fill_2
XFILLER_24_515 VPWR VGND sg13g2_fill_2
X_3926_ net705 _1034_ _1819_ VPWR VGND sg13g2_and2_1
X_3857_ _1775_ VPWR _0394_ VGND _1776_ _1777_ sg13g2_o21ai_1
X_2808_ _1049_ net825 _1043_ VPWR VGND sg13g2_xnor2_1
X_3788_ _1726_ _1720_ net862 _0933_ net428 VPWR VGND sg13g2_a22oi_1
XFILLER_30_1012 VPWR VGND sg13g2_decap_8
XFILLER_30_1023 VPWR VGND sg13g2_fill_2
X_2739_ _0987_ u_usb_cdc.u_sie.pid_q\[3\] _0986_ VPWR VGND sg13g2_xnor2_1
X_4409_ net727 VGND VPWR net853 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_2
XFILLER_46_128 VPWR VGND sg13g2_fill_2
XFILLER_28_832 VPWR VGND sg13g2_decap_4
XFILLER_42_312 VPWR VGND sg13g2_decap_8
XFILLER_15_559 VPWR VGND sg13g2_fill_1
XFILLER_24_74 VPWR VGND sg13g2_decap_4
XFILLER_7_747 VPWR VGND sg13g2_decap_8
XFILLER_10_297 VPWR VGND sg13g2_fill_2
XFILLER_3_920 VPWR VGND sg13g2_decap_8
XFILLER_2_441 VPWR VGND sg13g2_decap_8
XFILLER_3_997 VPWR VGND sg13g2_decap_8
XFILLER_38_607 VPWR VGND sg13g2_fill_1
XFILLER_19_843 VPWR VGND sg13g2_fill_1
XFILLER_18_375 VPWR VGND sg13g2_fill_1
XFILLER_18_386 VPWR VGND sg13g2_decap_4
XFILLER_33_334 VPWR VGND sg13g2_fill_1
XFILLER_34_868 VPWR VGND sg13g2_decap_4
XFILLER_33_367 VPWR VGND sg13g2_fill_1
XFILLER_14_570 VPWR VGND sg13g2_fill_2
X_3711_ _1529_ _1679_ _1680_ VPWR VGND sg13g2_nor2_1
X_3642_ VGND VPWR _1611_ _1613_ _1614_ net788 sg13g2_a21oi_1
X_3573_ VGND VPWR _1546_ _1547_ _1548_ net770 sg13g2_a21oi_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
XFILLER_5_290 VPWR VGND sg13g2_decap_8
X_2524_ VGND VPWR _0819_ _0683_ _0680_ sg13g2_or2_1
X_2455_ u_usb_cdc.u_ctrl_endp.req_q\[2\] u_usb_cdc.u_ctrl_endp.req_q\[8\] _0752_ VPWR
+ VGND sg13g2_nor2_2
X_2386_ _0550_ _0653_ net736 _0686_ VPWR VGND sg13g2_nand3_1
Xhold19 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[20\] VPWR VGND
+ net61 sg13g2_dlygate4sd3_1
X_4125_ net657 VGND VPWR net57 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[45\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_29_618 VPWR VGND sg13g2_fill_1
X_4056_ net731 VGND VPWR net353 _0051_ clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_43_109 VPWR VGND sg13g2_fill_2
X_3007_ _1147_ net104 _1146_ VPWR VGND sg13g2_nand2_1
X_3909_ net735 net234 _1804_ VPWR VGND sg13g2_nor2_1
XFILLER_4_739 VPWR VGND sg13g2_decap_8
XFILLER_3_205 VPWR VGND sg13g2_fill_1
XFILLER_0_934 VPWR VGND sg13g2_decap_8
XFILLER_48_938 VPWR VGND sg13g2_decap_8
XFILLER_19_52 VPWR VGND sg13g2_fill_1
XFILLER_16_835 VPWR VGND sg13g2_fill_1
XFILLER_34_109 VPWR VGND sg13g2_fill_1
XFILLER_16_868 VPWR VGND sg13g2_decap_8
XFILLER_31_816 VPWR VGND sg13g2_decap_4
XFILLER_24_890 VPWR VGND sg13g2_fill_2
XFILLER_31_838 VPWR VGND sg13g2_fill_2
XFILLER_35_95 VPWR VGND sg13g2_decap_8
XFILLER_3_794 VPWR VGND sg13g2_decap_8
X_2240_ _0542_ _1915_ VPWR VGND _0541_ sg13g2_nand2b_2
X_2171_ _0473_ u_usb_cdc.sie_out_data\[2\] net753 VPWR VGND sg13g2_xnor2_1
XFILLER_18_4 VPWR VGND sg13g2_fill_2
XFILLER_38_426 VPWR VGND sg13g2_fill_1
XFILLER_39_938 VPWR VGND sg13g2_decap_8
XFILLER_20_1022 VPWR VGND sg13g2_decap_8
XFILLER_47_982 VPWR VGND sg13g2_decap_8
XFILLER_21_348 VPWR VGND sg13g2_decap_8
X_3625_ net778 VPWR _1598_ VGND net786 net781 sg13g2_o21ai_1
X_3556_ _1487_ VPWR _0339_ VGND _1530_ _1531_ sg13g2_o21ai_1
X_2507_ _0714_ _0739_ _0803_ _0804_ VPWR VGND sg13g2_nor3_1
X_3487_ _0611_ net339 _1480_ VPWR VGND sg13g2_xor2_1
X_2438_ _0736_ net634 _0735_ VPWR VGND sg13g2_nand2_2
XFILLER_5_1027 VPWR VGND sg13g2_fill_2
XFILLER_5_1016 VPWR VGND sg13g2_decap_8
X_2369_ net770 net777 _0669_ VPWR VGND sg13g2_nor2b_1
XFILLER_45_919 VPWR VGND sg13g2_decap_8
X_4108_ net671 VGND VPWR net482 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[28\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
X_4039_ net678 VGND VPWR net872 u_usb_cdc.u_ctrl_endp.state_q\[3\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_2
XFILLER_25_665 VPWR VGND sg13g2_fill_2
XFILLER_40_624 VPWR VGND sg13g2_fill_2
XFILLER_13_827 VPWR VGND sg13g2_decap_8
XFILLER_40_646 VPWR VGND sg13g2_decap_4
XFILLER_21_64 VPWR VGND sg13g2_fill_1
XFILLER_21_97 VPWR VGND sg13g2_decap_8
XFILLER_0_731 VPWR VGND sg13g2_decap_8
XFILLER_48_735 VPWR VGND sg13g2_decap_8
XFILLER_47_212 VPWR VGND sg13g2_decap_4
XFILLER_36_908 VPWR VGND sg13g2_fill_2
XFILLER_47_289 VPWR VGND sg13g2_fill_1
XFILLER_29_993 VPWR VGND sg13g2_decap_8
XFILLER_44_941 VPWR VGND sg13g2_decap_8
XFILLER_31_613 VPWR VGND sg13g2_decap_8
XFILLER_31_646 VPWR VGND sg13g2_decap_4
XFILLER_8_842 VPWR VGND sg13g2_fill_2
XFILLER_7_330 VPWR VGND sg13g2_decap_4
XFILLER_12_893 VPWR VGND sg13g2_decap_8
Xhold308 _0337_ VPWR VGND net350 sg13g2_dlygate4sd3_1
XFILLER_8_875 VPWR VGND sg13g2_decap_8
XFILLER_7_352 VPWR VGND sg13g2_decap_8
X_4390_ net722 VGND VPWR _0392_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[11\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_2
Xhold319 _0419_ VPWR VGND net361 sg13g2_dlygate4sd3_1
X_3410_ _0548_ _0660_ _1429_ VPWR VGND sg13g2_nor2_1
X_3341_ net926 net392 _1384_ _0270_ VPWR VGND sg13g2_mux2_1
X_3272_ VGND VPWR net809 _1335_ _1338_ _1337_ sg13g2_a21oi_1
X_2223_ u_usb_cdc.u_sie.crc16_q\[3\] u_usb_cdc.u_sie.crc16_q\[2\] _0524_ _0525_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_39_735 VPWR VGND sg13g2_fill_2
X_2154_ _0457_ net635 _1958_ net703 net351 VPWR VGND sg13g2_a22oi_1
X_2085_ _1964_ net1069 VPWR VGND sg13g2_inv_2
XFILLER_35_985 VPWR VGND sg13g2_decap_8
X_2987_ _1135_ net709 _1134_ VPWR VGND sg13g2_nand2_2
X_3608_ _1559_ VPWR _0341_ VGND _1580_ _1581_ sg13g2_o21ai_1
X_3539_ VGND VPWR _0650_ _0661_ _1515_ _1440_ sg13g2_a21oi_1
XFILLER_27_1006 VPWR VGND sg13g2_decap_8
XFILLER_29_223 VPWR VGND sg13g2_decap_8
XFILLER_18_919 VPWR VGND sg13g2_fill_2
XFILLER_26_930 VPWR VGND sg13g2_fill_1
XFILLER_16_42 VPWR VGND sg13g2_fill_1
XFILLER_41_933 VPWR VGND sg13g2_decap_8
XFILLER_13_635 VPWR VGND sg13g2_fill_1
XFILLER_13_668 VPWR VGND sg13g2_fill_2
XFILLER_40_487 VPWR VGND sg13g2_fill_2
XFILLER_32_41 VPWR VGND sg13g2_fill_2
XFILLER_40_498 VPWR VGND sg13g2_decap_4
XFILLER_5_834 VPWR VGND sg13g2_decap_8
XFILLER_4_333 VPWR VGND sg13g2_decap_8
XFILLER_48_565 VPWR VGND sg13g2_decap_4
X_2910_ _1102_ net83 _1101_ VPWR VGND sg13g2_nand2_1
XFILLER_31_410 VPWR VGND sg13g2_decap_8
X_3890_ _1799_ VPWR _0405_ VGND _1937_ _0448_ sg13g2_o21ai_1
XFILLER_32_999 VPWR VGND sg13g2_decap_8
X_2841_ _1060_ VPWR _0091_ VGND _1062_ net616 sg13g2_o21ai_1
X_2772_ _1017_ _1016_ u_usb_cdc.u_sie.in_toggle_q\[2\] net633 u_usb_cdc.u_sie.in_toggle_q\[1\]
+ VPWR VGND sg13g2_a22oi_1
Xhold105 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[22\] VPWR VGND
+ net147 sg13g2_dlygate4sd3_1
Xhold116 _0171_ VPWR VGND net158 sg13g2_dlygate4sd3_1
XFILLER_7_193 VPWR VGND sg13g2_decap_4
X_4442_ net699 VGND VPWR net328 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
Xhold149 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[10\] VPWR VGND
+ net191 sg13g2_dlygate4sd3_1
Xhold138 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[14\] VPWR
+ VGND net180 sg13g2_dlygate4sd3_1
Xhold127 u_usb_cdc.u_sie.out_toggle_q\[0\] VPWR VGND net169 sg13g2_dlygate4sd3_1
X_4373_ net730 VGND VPWR _0375_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_2
Xfanout618 _0711_ net618 VPWR VGND sg13g2_buf_8
Xfanout629 _1220_ net629 VPWR VGND sg13g2_buf_8
Xfanout607 _1193_ net607 VPWR VGND sg13g2_buf_8
X_3324_ net619 _0662_ _1376_ VPWR VGND sg13g2_nor2_1
X_3255_ net805 net601 _1322_ _1323_ VPWR VGND sg13g2_nor3_1
XFILLER_39_510 VPWR VGND sg13g2_fill_2
X_2206_ _0508_ _0503_ _0506_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
X_3186_ _1261_ _0735_ _1242_ VPWR VGND sg13g2_nand2_1
X_2137_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\]
+ _0440_ VPWR VGND sg13g2_nor2_2
X_2068_ VPWR _1947_ net918 VGND sg13g2_inv_1
XFILLER_33_1021 VPWR VGND sg13g2_decap_8
Xhold672 _0261_ VPWR VGND net990 sg13g2_dlygate4sd3_1
XFILLER_2_837 VPWR VGND sg13g2_decap_8
Xhold650 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[1\] VPWR VGND
+ net968 sg13g2_dlygate4sd3_1
Xhold661 u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] VPWR VGND net979 sg13g2_dlygate4sd3_1
Xhold683 _1873_ VPWR VGND net1001 sg13g2_dlygate4sd3_1
XFILLER_1_358 VPWR VGND sg13g2_decap_8
Xhold694 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] VPWR VGND net1012 sg13g2_dlygate4sd3_1
XFILLER_17_204 VPWR VGND sg13g2_fill_1
XFILLER_17_226 VPWR VGND sg13g2_fill_2
XFILLER_14_988 VPWR VGND sg13g2_decap_8
XFILLER_13_487 VPWR VGND sg13g2_fill_2
XFILLER_49_830 VPWR VGND sg13g2_decap_8
X_3040_ VGND VPWR net611 _1170_ _0184_ _1169_ sg13g2_a21oi_1
XFILLER_36_557 VPWR VGND sg13g2_decap_8
X_3942_ _1827_ VPWR _0423_ VGND _1826_ _1833_ sg13g2_o21ai_1
X_3873_ _1788_ net704 net994 _0399_ VPWR VGND sg13g2_mux2_1
XFILLER_31_273 VPWR VGND sg13g2_decap_4
X_2824_ net9 net1039 net637 _0082_ VPWR VGND sg13g2_mux2_1
X_2755_ _1002_ net849 _1001_ VPWR VGND sg13g2_xnor2_1
X_2686_ _0951_ _0948_ net497 _1983_ net740 VPWR VGND sg13g2_a22oi_1
X_4425_ net725 VGND VPWR net44 u_usb_cdc.u_sie.u_phy_rx.dp_q\[1\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
X_4356_ net642 VGND VPWR net506 net17 clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3307_ _1358_ _1362_ _1363_ VPWR VGND sg13g2_nor2_1
X_4287_ net666 VGND VPWR _0289_ u_usb_cdc.u_ctrl_endp.max_length_q\[1\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_3238_ _1307_ net812 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[43\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_27_502 VPWR VGND sg13g2_decap_8
X_3169_ _1245_ net708 _1183_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_741 VPWR VGND sg13g2_fill_2
XFILLER_23_785 VPWR VGND sg13g2_fill_2
XFILLER_10_435 VPWR VGND sg13g2_fill_2
XFILLER_10_446 VPWR VGND sg13g2_fill_1
XFILLER_13_54 VPWR VGND sg13g2_decap_8
XFILLER_13_98 VPWR VGND sg13g2_decap_8
XFILLER_1_111 VPWR VGND sg13g2_fill_1
XFILLER_2_634 VPWR VGND sg13g2_decap_8
Xhold480 _0047_ VPWR VGND net522 sg13g2_dlygate4sd3_1
XFILLER_1_166 VPWR VGND sg13g2_fill_1
Xhold491 u_usb_cdc.out_valid_o[0] VPWR VGND net533 sg13g2_dlygate4sd3_1
XFILLER_49_126 VPWR VGND sg13g2_decap_8
XFILLER_1_199 VPWR VGND sg13g2_fill_2
XFILLER_46_844 VPWR VGND sg13g2_decap_8
XFILLER_45_332 VPWR VGND sg13g2_fill_2
XFILLER_33_516 VPWR VGND sg13g2_decap_8
XFILLER_14_752 VPWR VGND sg13g2_fill_2
XFILLER_6_940 VPWR VGND sg13g2_decap_8
X_2540_ _0833_ net845 _0832_ VPWR VGND sg13g2_nand2_1
XFILLER_5_472 VPWR VGND sg13g2_decap_8
X_2471_ VGND VPWR net760 _1926_ _0768_ _0710_ sg13g2_a21oi_1
X_4210_ net646 VGND VPWR net198 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[46\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4141_ net650 VGND VPWR net484 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[61\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_4072_ net648 VGND VPWR _0075_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_2
X_3023_ net823 _1150_ net754 _1159_ VPWR VGND sg13g2_nand3_1
XFILLER_24_538 VPWR VGND sg13g2_decap_8
X_3925_ _1818_ net705 _1034_ VPWR VGND sg13g2_nand2_2
XFILLER_20_733 VPWR VGND sg13g2_fill_1
X_3856_ net600 VPWR _1777_ VGND net366 _1773_ sg13g2_o21ai_1
X_2807_ _1047_ VPWR _1048_ VGND net707 _1043_ sg13g2_o21ai_1
XFILLER_20_799 VPWR VGND sg13g2_fill_1
X_3787_ VPWR _0376_ net429 VGND sg13g2_inv_1
XFILLER_3_409 VPWR VGND sg13g2_decap_8
X_2738_ VGND VPWR u_usb_cdc.endp\[0\] u_usb_cdc.u_sie.out_toggle_q\[1\] _0986_ _0985_
+ sg13g2_a21oi_1
X_4408_ net731 VGND VPWR net914 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_2
X_2669_ _0917_ _0937_ _0938_ VPWR VGND sg13g2_nor2_1
X_4339_ net685 VGND VPWR _0341_ u_usb_cdc.u_sie.data_q\[2\] clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_46_107 VPWR VGND sg13g2_decap_4
XFILLER_15_505 VPWR VGND sg13g2_decap_4
XFILLER_27_387 VPWR VGND sg13g2_fill_2
XFILLER_10_221 VPWR VGND sg13g2_fill_1
XFILLER_7_726 VPWR VGND sg13g2_decap_8
XFILLER_40_85 VPWR VGND sg13g2_fill_2
XFILLER_2_420 VPWR VGND sg13g2_decap_8
XFILLER_3_976 VPWR VGND sg13g2_decap_8
Xfanout790 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[2\] net790
+ VPWR VGND sg13g2_buf_8
XFILLER_18_321 VPWR VGND sg13g2_fill_2
XFILLER_18_332 VPWR VGND sg13g2_fill_2
XFILLER_19_866 VPWR VGND sg13g2_fill_2
XFILLER_19_877 VPWR VGND sg13g2_decap_8
XFILLER_34_836 VPWR VGND sg13g2_decap_4
X_3710_ _1679_ _1573_ u_usb_cdc.u_ctrl_endp.req_q\[2\] _1517_ _0672_ VPWR VGND sg13g2_a22oi_1
X_3641_ VGND VPWR net793 _1612_ _1613_ _1913_ sg13g2_a21oi_1
X_3572_ VGND VPWR _1543_ _1545_ _1547_ _0668_ sg13g2_a21oi_1
X_2523_ _0816_ VPWR _0006_ VGND _0802_ _0818_ sg13g2_o21ai_1
X_2454_ u_usb_cdc.u_ctrl_endp.req_q\[1\] _0747_ _0750_ _0751_ VPWR VGND sg13g2_nor3_1
X_2385_ _0685_ _0550_ _0653_ VPWR VGND sg13g2_nand2_1
XFILLER_39_0 VPWR VGND sg13g2_fill_1
X_4124_ net669 VGND VPWR net131 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[44\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_48_clk clknet_3_4__leaf_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
X_4055_ net694 VGND VPWR _0019_ u_usb_cdc.u_sie.phy_state_q\[11\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
X_3006_ net823 net709 net735 _1146_ VPWR VGND _1134_ sg13g2_nand4_1
XFILLER_37_663 VPWR VGND sg13g2_decap_8
XFILLER_25_869 VPWR VGND sg13g2_decap_8
XFILLER_24_346 VPWR VGND sg13g2_fill_2
XFILLER_33_880 VPWR VGND sg13g2_fill_2
XFILLER_20_541 VPWR VGND sg13g2_decap_4
X_3908_ VGND VPWR net360 net599 _0419_ _1803_ sg13g2_a21oi_1
X_3839_ _1764_ net710 net393 VPWR VGND sg13g2_nand2_1
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_10_33 VPWR VGND sg13g2_fill_1
XFILLER_0_913 VPWR VGND sg13g2_decap_8
XFILLER_48_917 VPWR VGND sg13g2_decap_8
XFILLER_19_86 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_39_clk clknet_3_5__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_27_140 VPWR VGND sg13g2_decap_8
XFILLER_43_622 VPWR VGND sg13g2_fill_2
XFILLER_35_41 VPWR VGND sg13g2_decap_8
XFILLER_11_552 VPWR VGND sg13g2_decap_4
XFILLER_7_545 VPWR VGND sg13g2_decap_8
XFILLER_3_773 VPWR VGND sg13g2_decap_8
XFILLER_2_261 VPWR VGND sg13g2_fill_1
XFILLER_39_917 VPWR VGND sg13g2_decap_8
X_2170_ _0472_ _0470_ _0471_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_961 VPWR VGND sg13g2_decap_8
XFILLER_19_663 VPWR VGND sg13g2_fill_1
XFILLER_19_674 VPWR VGND sg13g2_fill_2
XFILLER_22_839 VPWR VGND sg13g2_decap_8
XFILLER_33_176 VPWR VGND sg13g2_fill_2
X_3624_ VGND VPWR _1597_ _1596_ _1594_ sg13g2_or2_1
X_3555_ net597 VPWR _1531_ VGND net967 net624 sg13g2_o21ai_1
X_3486_ _1479_ net339 net594 VPWR VGND sg13g2_nand2_1
XFILLER_0_209 VPWR VGND sg13g2_decap_4
X_2506_ _1928_ _0726_ _0803_ VPWR VGND sg13g2_and2_1
X_2437_ net747 net750 _0604_ _0735_ VPWR VGND sg13g2_nor3_2
X_2368_ net774 _0667_ _0668_ VPWR VGND sg13g2_and2_1
X_4107_ net656 VGND VPWR net453 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[27\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2299_ net745 u_usb_cdc.u_sie.phy_state_q\[9\] _0601_ VPWR VGND sg13g2_nor2b_2
X_4038_ net678 VGND VPWR _0012_ u_usb_cdc.u_ctrl_endp.state_q\[2\] clknet_leaf_48_clk
+ sg13g2_dfrbpq_2
XFILLER_25_622 VPWR VGND sg13g2_decap_8
XFILLER_37_471 VPWR VGND sg13g2_decap_8
XFILLER_40_603 VPWR VGND sg13g2_fill_1
XFILLER_21_54 VPWR VGND sg13g2_fill_1
XFILLER_0_710 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_0_787 VPWR VGND sg13g2_decap_8
XFILLER_47_246 VPWR VGND sg13g2_decap_4
XFILLER_29_972 VPWR VGND sg13g2_decap_8
XFILLER_35_408 VPWR VGND sg13g2_fill_1
XFILLER_44_920 VPWR VGND sg13g2_decap_8
XFILLER_28_493 VPWR VGND sg13g2_fill_2
XFILLER_44_997 VPWR VGND sg13g2_decap_8
XFILLER_15_154 VPWR VGND sg13g2_fill_2
XFILLER_30_124 VPWR VGND sg13g2_decap_4
XFILLER_12_850 VPWR VGND sg13g2_fill_1
XFILLER_8_854 VPWR VGND sg13g2_decap_8
Xhold309 _0051_ VPWR VGND net351 sg13g2_dlygate4sd3_1
X_3340_ net880 net391 _1384_ _0269_ VPWR VGND sg13g2_mux2_1
X_3271_ net807 VPWR _1337_ VGND net810 _1334_ sg13g2_o21ai_1
XFILLER_30_4 VPWR VGND sg13g2_fill_2
X_2222_ _1951_ _1952_ _1950_ _0524_ VPWR VGND _1953_ sg13g2_nand4_1
X_2153_ VGND VPWR _2008_ _2011_ _0456_ net351 sg13g2_a21oi_1
XFILLER_27_909 VPWR VGND sg13g2_fill_1
XFILLER_38_213 VPWR VGND sg13g2_decap_4
XFILLER_26_419 VPWR VGND sg13g2_fill_2
XFILLER_19_482 VPWR VGND sg13g2_decap_4
XFILLER_19_493 VPWR VGND sg13g2_decap_4
X_2084_ _1963_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[2\]
+ VPWR VGND sg13g2_inv_2
XFILLER_34_430 VPWR VGND sg13g2_decap_8
XFILLER_35_964 VPWR VGND sg13g2_decap_8
XFILLER_34_463 VPWR VGND sg13g2_fill_1
X_2986_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\]
+ _1134_ VPWR VGND sg13g2_nor2_2
X_3607_ net597 VPWR _1581_ VGND net945 net624 sg13g2_o21ai_1
X_3538_ net777 _0549_ net780 _1514_ VPWR VGND sg13g2_nand3_1
X_3469_ net712 _1465_ _1468_ VPWR VGND sg13g2_nor2_1
XFILLER_29_257 VPWR VGND sg13g2_fill_2
XFILLER_44_238 VPWR VGND sg13g2_fill_2
XFILLER_41_912 VPWR VGND sg13g2_decap_8
XFILLER_25_463 VPWR VGND sg13g2_decap_8
XFILLER_41_989 VPWR VGND sg13g2_decap_8
XFILLER_5_813 VPWR VGND sg13g2_decap_8
XFILLER_48_544 VPWR VGND sg13g2_decap_8
XFILLER_0_584 VPWR VGND sg13g2_decap_8
X_2840_ net707 _1063_ net736 _1064_ VPWR VGND sg13g2_nand3_1
XFILLER_32_978 VPWR VGND sg13g2_decap_8
X_2771_ u_usb_cdc.endp\[0\] _1907_ u_usb_cdc.endp\[3\] u_usb_cdc.endp\[2\] _1016_
+ VPWR VGND sg13g2_nor4_1
Xhold106 _0105_ VPWR VGND net148 sg13g2_dlygate4sd3_1
Xhold117 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[51\] VPWR VGND
+ net159 sg13g2_dlygate4sd3_1
XFILLER_7_172 VPWR VGND sg13g2_decap_8
X_4441_ net724 VGND VPWR net245 u_usb_cdc.u_sie.u_phy_rx.se0_q clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
Xhold139 _0181_ VPWR VGND net181 sg13g2_dlygate4sd3_1
Xhold128 _0989_ VPWR VGND net170 sg13g2_dlygate4sd3_1
X_4372_ net729 VGND VPWR _0374_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[2\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_2
Xfanout608 net610 net608 VPWR VGND sg13g2_buf_8
Xfanout619 net620 net619 VPWR VGND sg13g2_buf_8
X_3323_ _1375_ net788 _1358_ _0262_ VPWR VGND sg13g2_mux2_1
X_3254_ VPWR VGND _1279_ _1321_ _1318_ net808 _1322_ _1317_ sg13g2_a221oi_1
X_2205_ _0503_ _0506_ _0507_ VPWR VGND sg13g2_nor2b_1
X_3185_ _1259_ VPWR _1260_ VGND net768 _1962_ sg13g2_o21ai_1
XFILLER_39_577 VPWR VGND sg13g2_fill_1
X_2136_ _2008_ _2009_ _2010_ _2012_ VGND VPWR _2011_ sg13g2_nor4_2
X_2067_ _1946_ net409 VPWR VGND sg13g2_inv_2
XFILLER_41_208 VPWR VGND sg13g2_fill_1
XFILLER_23_912 VPWR VGND sg13g2_decap_8
XFILLER_23_923 VPWR VGND sg13g2_fill_1
XFILLER_22_444 VPWR VGND sg13g2_fill_2
XFILLER_22_477 VPWR VGND sg13g2_fill_2
XFILLER_33_1000 VPWR VGND sg13g2_decap_8
X_2969_ net901 _1126_ _1123_ _0157_ VPWR VGND sg13g2_mux2_1
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_2_816 VPWR VGND sg13g2_decap_8
Xhold640 u_usb_cdc.endp\[1\] VPWR VGND net958 sg13g2_dlygate4sd3_1
Xhold651 _0252_ VPWR VGND net969 sg13g2_dlygate4sd3_1
Xhold662 u_usb_cdc.u_sie.data_q\[4\] VPWR VGND net980 sg13g2_dlygate4sd3_1
Xhold673 u_usb_cdc.sie_out_data\[6\] VPWR VGND net991 sg13g2_dlygate4sd3_1
Xhold684 u_usb_cdc.endp\[2\] VPWR VGND net1002 sg13g2_dlygate4sd3_1
Xhold695 _0030_ VPWR VGND net1013 sg13g2_dlygate4sd3_1
XFILLER_40_1026 VPWR VGND sg13g2_fill_2
XFILLER_18_706 VPWR VGND sg13g2_fill_1
XFILLER_18_739 VPWR VGND sg13g2_decap_8
XFILLER_14_967 VPWR VGND sg13g2_fill_2
XFILLER_13_477 VPWR VGND sg13g2_fill_2
XFILLER_14_978 VPWR VGND sg13g2_fill_1
XFILLER_0_381 VPWR VGND sg13g2_decap_8
XFILLER_49_886 VPWR VGND sg13g2_decap_8
XFILLER_36_503 VPWR VGND sg13g2_fill_2
XFILLER_16_260 VPWR VGND sg13g2_decap_8
X_3941_ _1832_ VPWR _1833_ VGND u_usb_cdc.u_sie.u_phy_tx.data_q\[3\] _1819_ sg13g2_o21ai_1
X_3872_ VGND VPWR _0934_ _1788_ _0937_ _0935_ sg13g2_a21oi_2
X_2823_ net8 net1042 net637 _0081_ VPWR VGND sg13g2_mux2_1
X_2754_ _0987_ _0998_ _0999_ _1000_ _1001_ VPWR VGND sg13g2_nor4_1
XFILLER_31_296 VPWR VGND sg13g2_decap_8
X_2685_ net343 VPWR _0033_ VGND _1960_ _0948_ sg13g2_o21ai_1
X_4424_ net727 VGND VPWR net47 u_usb_cdc.u_sie.u_phy_rx.dp_q\[0\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
X_4355_ net641 VGND VPWR net375 net16 clknet_leaf_4_clk sg13g2_dfrbpq_1
X_3306_ _1359_ VPWR _1362_ VGND net803 _1361_ sg13g2_o21ai_1
X_4286_ net666 VGND VPWR _0288_ u_usb_cdc.u_ctrl_endp.max_length_q\[0\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_3237_ net325 net164 net812 _1306_ VPWR VGND sg13g2_mux2_1
X_3168_ _1244_ net810 _1242_ VPWR VGND sg13g2_xnor2_1
X_2119_ VGND VPWR _1997_ _1995_ u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] sg13g2_or2_1
XFILLER_42_506 VPWR VGND sg13g2_decap_8
X_3099_ _1205_ net132 _1202_ VPWR VGND sg13g2_nand2_1
XFILLER_23_731 VPWR VGND sg13g2_fill_1
XFILLER_11_959 VPWR VGND sg13g2_decap_8
XFILLER_13_22 VPWR VGND sg13g2_fill_2
XFILLER_2_613 VPWR VGND sg13g2_decap_8
Xhold481 u_usb_cdc.u_ctrl_endp.max_length_q\[2\] VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold470 _0141_ VPWR VGND net512 sg13g2_dlygate4sd3_1
Xhold492 _0042_ VPWR VGND net534 sg13g2_dlygate4sd3_1
XFILLER_46_823 VPWR VGND sg13g2_decap_8
XFILLER_18_569 VPWR VGND sg13g2_fill_1
XFILLER_33_528 VPWR VGND sg13g2_decap_4
XFILLER_13_230 VPWR VGND sg13g2_decap_8
XFILLER_13_241 VPWR VGND sg13g2_fill_1
XFILLER_10_981 VPWR VGND sg13g2_decap_8
XFILLER_6_996 VPWR VGND sg13g2_decap_8
X_2470_ u_usb_cdc.u_ctrl_endp.rec_q\[0\] _1927_ _0703_ _0766_ _0767_ VPWR VGND sg13g2_nor4_1
X_4140_ net668 VGND VPWR net488 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[60\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_4071_ net672 VGND VPWR net543 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_49_683 VPWR VGND sg13g2_decap_8
X_3022_ _1158_ net153 _1146_ VPWR VGND sg13g2_nand2_1
XFILLER_24_517 VPWR VGND sg13g2_fill_1
X_3924_ _2003_ net702 _1817_ VPWR VGND sg13g2_nor2_1
XFILLER_20_712 VPWR VGND sg13g2_fill_2
X_3855_ net366 _1773_ _1776_ VPWR VGND sg13g2_and2_1
X_2806_ _1047_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] _1040_
+ VPWR VGND sg13g2_nand2b_1
X_3786_ _1725_ _1720_ net428 net579 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[4\]
+ VPWR VGND sg13g2_a22oi_1
X_2737_ net767 net169 _0985_ VPWR VGND sg13g2_nor2b_1
X_2668_ _0914_ _0936_ _0441_ _0937_ VPWR VGND sg13g2_nand3_1
X_4407_ net731 VGND VPWR net974 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[0\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_2
XFILLER_8_1015 VPWR VGND sg13g2_decap_8
X_2599_ u_usb_cdc.u_sie.addr_q\[4\] u_usb_cdc.addr\[4\] _0880_ VPWR VGND sg13g2_xor2_1
X_4338_ net685 VGND VPWR _0340_ u_usb_cdc.u_sie.data_q\[1\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_4269_ net679 VGND VPWR _0271_ u_usb_cdc.addr\[3\] clknet_leaf_43_clk sg13g2_dfrbpq_2
XFILLER_27_366 VPWR VGND sg13g2_fill_2
XFILLER_27_377 VPWR VGND sg13g2_fill_1
XFILLER_43_859 VPWR VGND sg13g2_decap_8
XFILLER_43_848 VPWR VGND sg13g2_decap_8
XFILLER_11_701 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_fill_2
XFILLER_3_955 VPWR VGND sg13g2_decap_8
XFILLER_2_476 VPWR VGND sg13g2_decap_8
XFILLER_2_498 VPWR VGND sg13g2_decap_4
XFILLER_1_14 VPWR VGND sg13g2_decap_8
Xfanout780 net782 net780 VPWR VGND sg13g2_buf_8
Xfanout791 net792 net791 VPWR VGND sg13g2_buf_8
XFILLER_14_1009 VPWR VGND sg13g2_decap_8
X_3640_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[52\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[60\]
+ net801 _1612_ VPWR VGND sg13g2_mux2_1
X_3571_ _1504_ VPWR _1546_ VGND net780 _0548_ sg13g2_o21ai_1
X_2522_ _0798_ _0817_ _0726_ _0818_ VPWR VGND sg13g2_nand3_1
XFILLER_6_793 VPWR VGND sg13g2_decap_8
XFILLER_46_2 VPWR VGND sg13g2_fill_1
X_2453_ VPWR _0750_ _0749_ VGND sg13g2_inv_1
X_2384_ net714 net588 net585 _0682_ _0684_ VPWR VGND sg13g2_or4_1
X_4123_ net655 VGND VPWR net150 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[43\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
X_4054_ net695 VGND VPWR _0018_ u_usb_cdc.u_sie.phy_state_q\[10\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
XFILLER_49_491 VPWR VGND sg13g2_decap_8
X_3005_ _1145_ VPWR _0174_ VGND net717 net613 sg13g2_o21ai_1
XFILLER_37_642 VPWR VGND sg13g2_fill_1
XFILLER_24_303 VPWR VGND sg13g2_fill_1
X_3907_ u_usb_cdc.u_sie.rx_data\[7\] net599 _1803_ VPWR VGND sg13g2_nor2_1
X_3838_ _1761_ VPWR _0389_ VGND _1762_ _1763_ sg13g2_o21ai_1
XFILLER_20_597 VPWR VGND sg13g2_decap_8
X_3769_ _1713_ _0601_ _0623_ VPWR VGND sg13g2_nand2_1
XFILLER_0_969 VPWR VGND sg13g2_decap_8
XFILLER_28_620 VPWR VGND sg13g2_fill_1
XFILLER_16_826 VPWR VGND sg13g2_decap_8
XFILLER_15_336 VPWR VGND sg13g2_fill_2
XFILLER_43_656 VPWR VGND sg13g2_decap_8
XFILLER_43_689 VPWR VGND sg13g2_decap_8
XFILLER_24_892 VPWR VGND sg13g2_fill_1
XFILLER_30_306 VPWR VGND sg13g2_decap_8
XFILLER_11_520 VPWR VGND sg13g2_fill_1
XFILLER_23_380 VPWR VGND sg13g2_decap_8
XFILLER_23_391 VPWR VGND sg13g2_fill_2
XFILLER_13_1020 VPWR VGND sg13g2_decap_8
XFILLER_3_752 VPWR VGND sg13g2_decap_8
XFILLER_32_8 VPWR VGND sg13g2_fill_1
XFILLER_47_940 VPWR VGND sg13g2_decap_8
XFILLER_18_6 VPWR VGND sg13g2_fill_1
XFILLER_21_317 VPWR VGND sg13g2_decap_8
X_3623_ _1595_ VPWR _1596_ VGND _0738_ _1593_ sg13g2_o21ai_1
X_3554_ VGND VPWR _1527_ _1528_ _1530_ _1501_ sg13g2_a21oi_1
X_3485_ _1476_ VPWR _0321_ VGND _0894_ _1478_ sg13g2_o21ai_1
X_2505_ _0802_ _0800_ _0730_ VPWR VGND sg13g2_nand2b_1
X_2436_ VGND VPWR _0734_ _0733_ net584 sg13g2_or2_1
X_2367_ net785 net783 _1915_ _0667_ VPWR VGND net778 sg13g2_nand4_1
X_4106_ net656 VGND VPWR net427 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[26\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2298_ _0600_ net832 net590 VPWR VGND sg13g2_nand2_1
X_4037_ net678 VGND VPWR net551 u_usb_cdc.u_ctrl_endp.state_q\[1\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
XFILLER_37_450 VPWR VGND sg13g2_fill_1
XFILLER_38_984 VPWR VGND sg13g2_decap_8
XFILLER_25_689 VPWR VGND sg13g2_fill_1
XFILLER_21_895 VPWR VGND sg13g2_fill_2
XFILLER_43_1013 VPWR VGND sg13g2_decap_8
XFILLER_0_766 VPWR VGND sg13g2_decap_8
XFILLER_46_85 VPWR VGND sg13g2_fill_2
XFILLER_44_976 VPWR VGND sg13g2_decap_8
XFILLER_43_486 VPWR VGND sg13g2_fill_2
XFILLER_31_659 VPWR VGND sg13g2_fill_1
XFILLER_8_822 VPWR VGND sg13g2_decap_4
X_3270_ VGND VPWR _1336_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[6\]
+ net813 sg13g2_or2_1
X_2221_ _0523_ _0502_ _0509_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_593 VPWR VGND sg13g2_decap_4
X_2152_ _0455_ _2008_ _2011_ VPWR VGND sg13g2_nand2_1
XFILLER_39_737 VPWR VGND sg13g2_fill_1
X_2083_ VPWR _1962_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\]
+ VGND sg13g2_inv_1
XFILLER_35_943 VPWR VGND sg13g2_decap_8
X_2985_ _1133_ VPWR _0166_ VGND _1914_ _1130_ sg13g2_o21ai_1
X_3606_ VPWR VGND _1528_ _1489_ _1579_ net631 _1580_ _1568_ sg13g2_a221oi_1
X_3537_ _0544_ VPWR _1513_ VGND _1510_ _1512_ sg13g2_o21ai_1
XFILLER_1_519 VPWR VGND sg13g2_decap_8
X_3468_ net742 _1466_ net1005 _1467_ VPWR VGND sg13g2_nand3_1
X_3399_ net890 net568 _1420_ VPWR VGND sg13g2_nor2_1
X_2419_ net714 net586 net584 _0701_ _0717_ VPWR VGND sg13g2_or4_1
XFILLER_29_247 VPWR VGND sg13g2_fill_2
XFILLER_45_729 VPWR VGND sg13g2_decap_8
XFILLER_44_228 VPWR VGND sg13g2_fill_1
XFILLER_44_217 VPWR VGND sg13g2_fill_2
XFILLER_16_11 VPWR VGND sg13g2_decap_4
XFILLER_16_33 VPWR VGND sg13g2_fill_1
XFILLER_13_604 VPWR VGND sg13g2_decap_8
XFILLER_26_987 VPWR VGND sg13g2_decap_8
XFILLER_41_968 VPWR VGND sg13g2_decap_8
XFILLER_40_423 VPWR VGND sg13g2_decap_8
XFILLER_40_434 VPWR VGND sg13g2_fill_1
XFILLER_8_129 VPWR VGND sg13g2_fill_2
XFILLER_10_1023 VPWR VGND sg13g2_decap_4
XFILLER_5_869 VPWR VGND sg13g2_decap_8
XFILLER_0_563 VPWR VGND sg13g2_decap_8
XFILLER_48_523 VPWR VGND sg13g2_decap_8
XFILLER_16_442 VPWR VGND sg13g2_decap_8
XFILLER_28_280 VPWR VGND sg13g2_fill_2
XFILLER_16_475 VPWR VGND sg13g2_decap_4
XFILLER_32_957 VPWR VGND sg13g2_decap_8
XFILLER_31_445 VPWR VGND sg13g2_fill_2
X_2770_ _1015_ net633 _1014_ VPWR VGND sg13g2_nand2_1
Xhold107 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[43\] VPWR VGND
+ net149 sg13g2_dlygate4sd3_1
X_4440_ net698 VGND VPWR _0431_ _0060_ clknet_leaf_30_clk sg13g2_dfrbpq_2
Xhold118 _0134_ VPWR VGND net160 sg13g2_dlygate4sd3_1
Xhold129 _0067_ VPWR VGND net171 sg13g2_dlygate4sd3_1
X_4371_ net728 VGND VPWR _0373_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[1\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
Xfanout609 net610 net609 VPWR VGND sg13g2_buf_1
X_3322_ _1373_ VPWR _1375_ VGND _1361_ _1374_ sg13g2_o21ai_1
X_3253_ _1278_ _1319_ _1320_ _1321_ VPWR VGND sg13g2_nor3_1
X_2204_ _0506_ _0504_ _0505_ VPWR VGND sg13g2_xnor2_1
X_3184_ _1259_ net768 net968 VPWR VGND sg13g2_nand2_1
XFILLER_14_0 VPWR VGND sg13g2_fill_1
X_2135_ _1935_ net913 _2011_ VPWR VGND sg13g2_nor2_1
XFILLER_27_729 VPWR VGND sg13g2_fill_2
X_2066_ VPWR _1945_ net881 VGND sg13g2_inv_1
XFILLER_23_902 VPWR VGND sg13g2_fill_1
XFILLER_22_423 VPWR VGND sg13g2_fill_1
X_2968_ _1052_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] _1054_
+ _1126_ VPWR VGND sg13g2_mux2_1
X_2899_ _1099_ net824 _1057_ VPWR VGND sg13g2_nand2_2
Xhold630 _0014_ VPWR VGND net948 sg13g2_dlygate4sd3_1
Xhold652 u_usb_cdc.u_ctrl_endp.req_q\[2\] VPWR VGND net970 sg13g2_dlygate4sd3_1
Xhold641 _0304_ VPWR VGND net959 sg13g2_dlygate4sd3_1
Xhold663 u_usb_cdc.u_sie.phy_state_q\[9\] VPWR VGND net981 sg13g2_dlygate4sd3_1
Xhold696 u_usb_cdc.sie_out_data\[5\] VPWR VGND net1014 sg13g2_dlygate4sd3_1
Xhold685 u_usb_cdc.u_ctrl_endp.state_q\[6\] VPWR VGND net1003 sg13g2_dlygate4sd3_1
Xhold674 u_usb_cdc.u_sie.rx_data\[5\] VPWR VGND net992 sg13g2_dlygate4sd3_1
XFILLER_40_1005 VPWR VGND sg13g2_decap_8
XFILLER_26_740 VPWR VGND sg13g2_decap_8
XFILLER_43_31 VPWR VGND sg13g2_fill_2
XFILLER_41_798 VPWR VGND sg13g2_decap_8
XFILLER_4_143 VPWR VGND sg13g2_fill_2
XFILLER_0_360 VPWR VGND sg13g2_decap_8
XFILLER_1_883 VPWR VGND sg13g2_decap_8
XFILLER_49_865 VPWR VGND sg13g2_decap_8
XFILLER_36_515 VPWR VGND sg13g2_fill_1
X_3940_ _1819_ VPWR _1832_ VGND net702 _1831_ sg13g2_o21ai_1
XFILLER_16_283 VPWR VGND sg13g2_fill_2
X_3871_ _0398_ _1787_ _1959_ _1786_ _0947_ VPWR VGND sg13g2_a22oi_1
XFILLER_31_242 VPWR VGND sg13g2_fill_1
XFILLER_32_776 VPWR VGND sg13g2_fill_2
X_2822_ net7 net1041 net637 _0080_ VPWR VGND sg13g2_mux2_1
X_2753_ _1000_ net633 net769 VPWR VGND sg13g2_nand2b_1
XFILLER_9_994 VPWR VGND sg13g2_decap_8
XFILLER_8_493 VPWR VGND sg13g2_decap_4
X_2684_ _0950_ net342 _0949_ VPWR VGND sg13g2_nand2_1
X_4423_ net734 VGND VPWR net236 u_usb_cdc.dp_pu_o clknet_leaf_4_clk sg13g2_dfrbpq_1
X_4354_ net641 VGND VPWR net421 net15 clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3305_ net631 u_usb_cdc.sie_in_req net626 _1361_ VPWR VGND sg13g2_a21o_1
X_4285_ net677 VGND VPWR _0287_ u_usb_cdc.u_ctrl_endp.in_dir_q clknet_leaf_50_clk
+ sg13g2_dfrbpq_2
X_3236_ _0245_ _1305_ _1304_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_353 VPWR VGND sg13g2_fill_2
X_3167_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\] _1183_
+ net820 _1243_ VPWR VGND sg13g2_nand3_1
XFILLER_39_364 VPWR VGND sg13g2_decap_4
X_3098_ _1204_ VPWR _0208_ VGND net708 _1153_ sg13g2_o21ai_1
X_2118_ u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] _1995_ _1996_ VPWR VGND sg13g2_nor2_1
X_2049_ VPWR _1928_ u_usb_cdc.u_ctrl_endp.in_dir_q VGND sg13g2_inv_1
XFILLER_23_776 VPWR VGND sg13g2_decap_4
XFILLER_11_938 VPWR VGND sg13g2_decap_8
XFILLER_22_275 VPWR VGND sg13g2_decap_8
XFILLER_10_437 VPWR VGND sg13g2_fill_1
Xhold460 u_usb_cdc.u_sie.crc16_q\[2\] VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold471 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[37\] VPWR VGND
+ net513 sg13g2_dlygate4sd3_1
XFILLER_2_669 VPWR VGND sg13g2_decap_8
Xhold482 _0290_ VPWR VGND net524 sg13g2_dlygate4sd3_1
Xhold493 _0049_ VPWR VGND net535 sg13g2_dlygate4sd3_1
XFILLER_46_802 VPWR VGND sg13g2_decap_8
XFILLER_45_345 VPWR VGND sg13g2_decap_4
XFILLER_45_334 VPWR VGND sg13g2_fill_1
XFILLER_46_879 VPWR VGND sg13g2_decap_8
XFILLER_14_710 VPWR VGND sg13g2_decap_8
XFILLER_14_721 VPWR VGND sg13g2_fill_1
XFILLER_14_754 VPWR VGND sg13g2_fill_1
XFILLER_9_268 VPWR VGND sg13g2_fill_1
XFILLER_9_279 VPWR VGND sg13g2_decap_4
XFILLER_10_960 VPWR VGND sg13g2_decap_8
XFILLER_6_975 VPWR VGND sg13g2_decap_8
XFILLER_1_680 VPWR VGND sg13g2_decap_8
X_4070_ net699 VGND VPWR net309 _0054_ clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_49_662 VPWR VGND sg13g2_decap_8
X_3021_ _1156_ VPWR _0178_ VGND net821 _1157_ sg13g2_o21ai_1
X_3923_ _1816_ net282 net621 VPWR VGND sg13g2_nand2_1
X_3854_ _1775_ net710 net366 VPWR VGND sg13g2_nand2_1
X_2805_ _1046_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[1\] _1045_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_20_768 VPWR VGND sg13g2_decap_8
X_3785_ VPWR _0375_ net528 VGND sg13g2_inv_1
X_2736_ VPWR _0984_ _0983_ VGND sg13g2_inv_1
X_2667_ _0442_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] _0936_ VPWR VGND sg13g2_nor2b_1
X_4406_ net728 VGND VPWR _0044_ u_usb_cdc.u_sie.u_phy_rx.rx_err_q clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_2598_ _0879_ u_usb_cdc.addr\[6\] net250 VPWR VGND sg13g2_xnor2_1
X_4337_ net685 VGND VPWR _0339_ u_usb_cdc.u_sie.data_q\[0\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_4268_ net693 VGND VPWR _0270_ u_usb_cdc.addr\[2\] clknet_leaf_43_clk sg13g2_dfrbpq_2
X_3219_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[1\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[9\]
+ net816 _1290_ VPWR VGND sg13g2_mux2_1
X_4199_ net644 VGND VPWR _0202_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[35\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_28_846 VPWR VGND sg13g2_fill_2
XFILLER_43_827 VPWR VGND sg13g2_decap_8
XFILLER_15_518 VPWR VGND sg13g2_fill_2
XFILLER_42_348 VPWR VGND sg13g2_fill_1
XFILLER_10_245 VPWR VGND sg13g2_fill_2
XFILLER_40_87 VPWR VGND sg13g2_fill_1
XFILLER_3_934 VPWR VGND sg13g2_decap_8
XFILLER_2_455 VPWR VGND sg13g2_decap_8
Xhold290 _0382_ VPWR VGND net332 sg13g2_dlygate4sd3_1
XFILLER_1_37 VPWR VGND sg13g2_fill_2
Xfanout770 net772 net770 VPWR VGND sg13g2_buf_8
Xfanout781 net782 net781 VPWR VGND sg13g2_buf_1
Xfanout792 net793 net792 VPWR VGND sg13g2_buf_8
XFILLER_46_698 VPWR VGND sg13g2_fill_2
XFILLER_42_893 VPWR VGND sg13g2_decap_8
XFILLER_41_381 VPWR VGND sg13g2_fill_2
XFILLER_10_790 VPWR VGND sg13g2_fill_1
X_3570_ VGND VPWR _1545_ _1544_ _1542_ sg13g2_or2_1
X_2521_ net884 net860 _0734_ _0736_ _0817_ VPWR VGND sg13g2_nor4_1
XFILLER_6_772 VPWR VGND sg13g2_decap_8
X_2452_ u_usb_cdc.u_ctrl_endp.req_q\[6\] net842 u_usb_cdc.u_ctrl_endp.req_q\[7\] _0749_
+ VPWR VGND sg13g2_nor3_1
X_2383_ net585 _0682_ _0683_ VPWR VGND sg13g2_nor2_1
X_4122_ net655 VGND VPWR net111 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[42\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_4053_ net694 VGND VPWR _0028_ u_usb_cdc.u_sie.phy_state_q\[9\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_49_470 VPWR VGND sg13g2_decap_8
X_3004_ _1145_ net229 net613 VPWR VGND sg13g2_nand2_1
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
XFILLER_25_827 VPWR VGND sg13g2_decap_8
XFILLER_25_838 VPWR VGND sg13g2_fill_2
X_3906_ net982 net908 net599 _0418_ VPWR VGND sg13g2_mux2_1
XFILLER_33_882 VPWR VGND sg13g2_fill_1
X_3837_ net600 VPWR _1763_ VGND net402 _1758_ sg13g2_o21ai_1
XFILLER_20_554 VPWR VGND sg13g2_fill_2
X_3768_ _1711_ net750 _1712_ _0370_ VPWR VGND sg13g2_a21o_1
X_2719_ net743 _0973_ _0045_ VPWR VGND sg13g2_nor2_1
X_3699_ _1667_ VPWR _1668_ VGND net801 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[7\]
+ sg13g2_o21ai_1
XFILLER_0_948 VPWR VGND sg13g2_decap_8
XFILLER_28_643 VPWR VGND sg13g2_decap_8
XFILLER_43_624 VPWR VGND sg13g2_fill_1
XFILLER_27_186 VPWR VGND sg13g2_decap_4
XFILLER_11_576 VPWR VGND sg13g2_fill_2
XFILLER_3_731 VPWR VGND sg13g2_decap_8
XFILLER_25_8 VPWR VGND sg13g2_decap_8
XFILLER_46_451 VPWR VGND sg13g2_fill_1
XFILLER_19_676 VPWR VGND sg13g2_fill_1
XFILLER_47_996 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_4
XFILLER_33_178 VPWR VGND sg13g2_fill_1
XFILLER_30_830 VPWR VGND sg13g2_decap_8
XFILLER_30_852 VPWR VGND sg13g2_fill_2
X_3622_ _0544_ u_usb_cdc.u_ctrl_endp.req_q\[8\] _1595_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_580 VPWR VGND sg13g2_fill_1
X_3553_ _0560_ _0576_ _0554_ _1529_ VPWR VGND sg13g2_nand3_1
X_3484_ _1478_ _0611_ _1477_ VPWR VGND sg13g2_nand2_1
XFILLER_44_0 VPWR VGND sg13g2_fill_1
X_2504_ _0801_ _0800_ _0788_ VPWR VGND sg13g2_nand2b_1
X_2435_ _0733_ u_usb_cdc.u_ctrl_endp.state_q\[2\] _0624_ VPWR VGND sg13g2_nand2_1
X_2366_ net773 _0665_ _0666_ VPWR VGND sg13g2_nor2_1
X_4105_ net653 VGND VPWR net490 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[25\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2297_ _1903_ _0528_ _0599_ VPWR VGND sg13g2_nor2_1
X_4036_ net678 VGND VPWR net537 _0049_ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_38_963 VPWR VGND sg13g2_decap_8
XFILLER_24_101 VPWR VGND sg13g2_fill_2
XFILLER_25_679 VPWR VGND sg13g2_fill_2
XFILLER_36_1010 VPWR VGND sg13g2_decap_8
XFILLER_20_362 VPWR VGND sg13g2_decap_8
XFILLER_0_745 VPWR VGND sg13g2_decap_8
XFILLER_48_749 VPWR VGND sg13g2_decap_8
XFILLER_28_440 VPWR VGND sg13g2_fill_2
XFILLER_44_955 VPWR VGND sg13g2_decap_8
XFILLER_15_156 VPWR VGND sg13g2_fill_1
XFILLER_24_690 VPWR VGND sg13g2_fill_1
XFILLER_11_362 VPWR VGND sg13g2_fill_2
XFILLER_12_885 VPWR VGND sg13g2_fill_2
XFILLER_8_889 VPWR VGND sg13g2_decap_8
XFILLER_3_572 VPWR VGND sg13g2_decap_8
X_2220_ VPWR _0522_ _0521_ VGND sg13g2_inv_1
XFILLER_30_6 VPWR VGND sg13g2_fill_1
XFILLER_16_4 VPWR VGND sg13g2_decap_8
X_2151_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] _1935_ net257 net635 _0454_ VPWR VGND
+ sg13g2_and4_1
X_2082_ VPWR _1961_ net987 VGND sg13g2_inv_1
XFILLER_47_793 VPWR VGND sg13g2_decap_8
XFILLER_35_999 VPWR VGND sg13g2_decap_8
XFILLER_21_104 VPWR VGND sg13g2_fill_2
X_2984_ _1133_ net335 _1130_ VPWR VGND sg13g2_nand2_1
XFILLER_30_660 VPWR VGND sg13g2_fill_2
X_3605_ _1574_ _1578_ _1579_ VPWR VGND sg13g2_nor2_1
X_3536_ VGND VPWR _0547_ _1511_ _1512_ net777 sg13g2_a21oi_1
X_3467_ net507 net1005 net460 _1466_ VPWR VGND _1465_ sg13g2_nand4_1
X_2418_ _0656_ net574 net715 _0716_ VPWR VGND net617 sg13g2_nand4_1
X_3398_ VGND VPWR net568 _1419_ _0293_ _1418_ sg13g2_a21oi_1
X_2349_ _0649_ _1917_ _0552_ VPWR VGND sg13g2_nand2_2
XFILLER_45_708 VPWR VGND sg13g2_decap_8
XFILLER_29_259 VPWR VGND sg13g2_fill_1
XFILLER_44_207 VPWR VGND sg13g2_fill_1
X_4019_ net686 VGND VPWR net171 u_usb_cdc.u_sie.out_toggle_q\[0\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_38_793 VPWR VGND sg13g2_fill_2
XFILLER_40_402 VPWR VGND sg13g2_fill_1
XFILLER_41_947 VPWR VGND sg13g2_decap_8
XFILLER_9_609 VPWR VGND sg13g2_decap_4
XFILLER_21_682 VPWR VGND sg13g2_decap_8
XFILLER_20_181 VPWR VGND sg13g2_fill_2
XFILLER_5_848 VPWR VGND sg13g2_decap_8
XFILLER_10_1002 VPWR VGND sg13g2_decap_8
XFILLER_48_502 VPWR VGND sg13g2_decap_8
XFILLER_0_542 VPWR VGND sg13g2_decap_8
XFILLER_29_771 VPWR VGND sg13g2_fill_2
XFILLER_31_424 VPWR VGND sg13g2_fill_2
XFILLER_40_991 VPWR VGND sg13g2_decap_8
XFILLER_12_671 VPWR VGND sg13g2_fill_1
XFILLER_8_653 VPWR VGND sg13g2_fill_1
Xhold108 _0126_ VPWR VGND net150 sg13g2_dlygate4sd3_1
Xhold119 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[63\] VPWR
+ VGND net161 sg13g2_dlygate4sd3_1
X_4370_ net728 VGND VPWR _0372_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
X_3321_ _1374_ _1914_ _1368_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_391 VPWR VGND sg13g2_fill_1
X_3252_ net816 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[20\]
+ _1320_ VPWR VGND sg13g2_nor2_1
X_2203_ net762 net563 _0505_ VPWR VGND sg13g2_xor2_1
X_3183_ net578 net822 _1258_ _0239_ VPWR VGND sg13g2_a21o_1
X_2134_ _1934_ net973 _2010_ VPWR VGND sg13g2_nor2_1
X_2065_ VPWR _1944_ net540 VGND sg13g2_inv_1
XFILLER_22_402 VPWR VGND sg13g2_decap_8
XFILLER_23_947 VPWR VGND sg13g2_fill_2
XFILLER_22_446 VPWR VGND sg13g2_fill_1
X_2967_ net857 _1125_ _1123_ _0156_ VPWR VGND sg13g2_mux2_1
X_2898_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ net473 _1098_ _0114_ VPWR VGND sg13g2_mux2_1
Xhold620 _0313_ VPWR VGND net938 sg13g2_dlygate4sd3_1
Xhold631 u_usb_cdc.u_ctrl_endp.req_q\[9\] VPWR VGND net949 sg13g2_dlygate4sd3_1
Xhold653 u_usb_cdc.u_ctrl_endp.req_q\[4\] VPWR VGND net971 sg13g2_dlygate4sd3_1
Xhold642 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[3\] VPWR VGND
+ net960 sg13g2_dlygate4sd3_1
Xhold675 u_usb_cdc.u_ctrl_endp.in_dir_q VPWR VGND net993 sg13g2_dlygate4sd3_1
Xhold697 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\] VPWR
+ VGND net1015 sg13g2_dlygate4sd3_1
Xhold686 _0016_ VPWR VGND net1004 sg13g2_dlygate4sd3_1
Xhold664 u_usb_cdc.u_sie.rx_data\[6\] VPWR VGND net982 sg13g2_dlygate4sd3_1
X_3519_ VGND VPWR net799 _1967_ _1495_ net792 sg13g2_a21oi_1
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
XFILLER_26_774 VPWR VGND sg13g2_fill_2
XFILLER_13_402 VPWR VGND sg13g2_decap_8
XFILLER_40_210 VPWR VGND sg13g2_fill_2
XFILLER_41_766 VPWR VGND sg13g2_fill_1
XFILLER_14_969 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_20_clk clknet_3_3__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_5_645 VPWR VGND sg13g2_fill_2
XFILLER_4_122 VPWR VGND sg13g2_fill_1
XFILLER_1_862 VPWR VGND sg13g2_decap_8
XFILLER_49_844 VPWR VGND sg13g2_decap_8
XFILLER_36_505 VPWR VGND sg13g2_fill_1
X_3870_ net600 _1782_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] _1787_ VPWR VGND sg13g2_nand3_1
XFILLER_17_1008 VPWR VGND sg13g2_decap_8
X_2821_ net6 net1033 net637 _0079_ VPWR VGND sg13g2_mux2_1
X_2752_ _0999_ _0594_ _0604_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_11_clk clknet_3_2__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_9_973 VPWR VGND sg13g2_decap_8
X_2683_ net393 net402 net740 _0949_ VPWR VGND sg13g2_nand3_1
X_4422_ net725 VGND VPWR net522 u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[1\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
X_4353_ net641 VGND VPWR _0355_ net14 clknet_leaf_4_clk sg13g2_dfrbpq_1
X_4284_ net666 VGND VPWR net885 u_usb_cdc.u_ctrl_endp.class_q clknet_leaf_50_clk sg13g2_dfrbpq_2
X_3304_ net803 net794 net790 _1914_ _1360_ VPWR VGND sg13g2_nor4_1
X_3235_ _1305_ _1296_ net120 net601 net495 VPWR VGND sg13g2_a22oi_1
XFILLER_39_310 VPWR VGND sg13g2_fill_1
X_3166_ net1015 net822 _1242_ VPWR VGND sg13g2_xor2_1
X_3097_ _1204_ net246 _1202_ VPWR VGND sg13g2_nand2_1
X_2117_ _1995_ u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[1\] u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[2\]
+ VPWR VGND sg13g2_nand2_1
X_2048_ _1927_ net910 VPWR VGND sg13g2_inv_2
XFILLER_11_917 VPWR VGND sg13g2_decap_8
XFILLER_13_24 VPWR VGND sg13g2_fill_1
X_3999_ _1880_ u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] net316 VPWR VGND sg13g2_xnor2_1
XFILLER_6_409 VPWR VGND sg13g2_decap_8
Xhold472 _0120_ VPWR VGND net514 sg13g2_dlygate4sd3_1
XFILLER_2_648 VPWR VGND sg13g2_decap_8
Xhold461 net20 VPWR VGND net503 sg13g2_dlygate4sd3_1
Xhold450 _0154_ VPWR VGND net492 sg13g2_dlygate4sd3_1
Xhold494 _0642_ VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold483 u_usb_cdc.u_sie.phy_state_q\[3\] VPWR VGND net525 sg13g2_dlygate4sd3_1
XFILLER_38_32 VPWR VGND sg13g2_fill_1
XFILLER_46_858 VPWR VGND sg13g2_decap_8
XFILLER_13_254 VPWR VGND sg13g2_decap_8
XFILLER_6_954 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_486 VPWR VGND sg13g2_fill_1
X_3020_ net823 _1150_ net755 _1157_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_36_357 VPWR VGND sg13g2_fill_1
XFILLER_45_891 VPWR VGND sg13g2_decap_8
X_3922_ _0421_ _1813_ _1815_ net622 _1975_ VPWR VGND sg13g2_a22oi_1
X_3853_ net887 net710 _1774_ _0393_ VPWR VGND sg13g2_a21o_1
X_2804_ net1053 net997 _1045_ VPWR VGND sg13g2_xor2_1
XFILLER_32_596 VPWR VGND sg13g2_decap_4
X_3784_ _1724_ _1720_ net527 net579 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_30_1005 VPWR VGND sg13g2_decap_8
XFILLER_8_291 VPWR VGND sg13g2_fill_1
X_2735_ _0980_ _0982_ _0983_ VPWR VGND sg13g2_and2_1
X_2666_ _0935_ net515 _0447_ VPWR VGND sg13g2_nand2_1
X_4405_ net729 VGND VPWR net978 u_usb_cdc.u_sie.rx_valid clknet_leaf_33_clk sg13g2_dfrbpq_1
X_4336_ net695 VGND VPWR _0338_ u_usb_cdc.u_sie.crc16_q\[15\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_2597_ u_usb_cdc.u_sie.addr_q\[0\] u_usb_cdc.addr\[0\] _0878_ VPWR VGND sg13g2_xor2_1
X_4267_ net680 VGND VPWR _0269_ u_usb_cdc.addr\[1\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_3218_ net815 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[33\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[41\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[49\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[57\] net811 _1289_
+ VPWR VGND sg13g2_mux4_1
X_4198_ net659 VGND VPWR _0201_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[34\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_28_803 VPWR VGND sg13g2_fill_1
X_3149_ _1232_ net145 _1230_ VPWR VGND sg13g2_nand2_1
XFILLER_28_836 VPWR VGND sg13g2_fill_1
XFILLER_23_541 VPWR VGND sg13g2_fill_2
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_24_78 VPWR VGND sg13g2_fill_1
XFILLER_6_206 VPWR VGND sg13g2_decap_4
XFILLER_11_769 VPWR VGND sg13g2_fill_1
XFILLER_40_44 VPWR VGND sg13g2_fill_1
XFILLER_3_913 VPWR VGND sg13g2_decap_8
XFILLER_46_1012 VPWR VGND sg13g2_decap_8
Xhold280 _0185_ VPWR VGND net322 sg13g2_dlygate4sd3_1
XFILLER_2_434 VPWR VGND sg13g2_decap_8
XFILLER_49_64 VPWR VGND sg13g2_decap_4
XFILLER_49_53 VPWR VGND sg13g2_decap_4
Xhold291 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[2\] VPWR VGND net333 sg13g2_dlygate4sd3_1
Xfanout760 net761 net760 VPWR VGND sg13g2_buf_8
Xfanout782 net783 net782 VPWR VGND sg13g2_buf_2
Xfanout771 net772 net771 VPWR VGND sg13g2_buf_1
Xfanout793 net796 net793 VPWR VGND sg13g2_buf_8
XFILLER_46_633 VPWR VGND sg13g2_fill_2
XFILLER_33_305 VPWR VGND sg13g2_decap_4
XFILLER_33_327 VPWR VGND sg13g2_decap_8
XFILLER_14_530 VPWR VGND sg13g2_decap_8
XFILLER_14_541 VPWR VGND sg13g2_fill_2
XFILLER_41_393 VPWR VGND sg13g2_fill_2
XFILLER_6_751 VPWR VGND sg13g2_decap_8
X_2520_ net842 VPWR _0816_ VGND _0720_ _0815_ sg13g2_o21ai_1
X_2451_ u_usb_cdc.u_ctrl_endp.req_q\[6\] net842 _0748_ VPWR VGND sg13g2_nor2_1
X_2382_ net841 u_usb_cdc.u_ctrl_endp.state_q\[6\] _0557_ _0681_ _0682_ VPWR VGND sg13g2_or4_1
X_4121_ net655 VGND VPWR net74 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[41\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4052_ net697 VGND VPWR net848 u_usb_cdc.u_sie.phy_state_q\[8\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_2
XFILLER_37_600 VPWR VGND sg13g2_fill_1
X_3003_ _1144_ VPWR _0173_ VGND _1901_ net614 sg13g2_o21ai_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
XFILLER_37_677 VPWR VGND sg13g2_decap_4
XFILLER_24_327 VPWR VGND sg13g2_decap_4
X_3905_ net992 net862 _0972_ _0417_ VPWR VGND sg13g2_mux2_1
X_3836_ net402 _1758_ _1762_ VPWR VGND sg13g2_and2_1
X_3767_ _1465_ _1708_ _1711_ _1712_ VPWR VGND sg13g2_nor3_1
X_2718_ net529 net599 _0973_ VPWR VGND sg13g2_nor2_1
X_3698_ VGND VPWR net801 _1973_ _1667_ net793 sg13g2_a21oi_1
X_2649_ _0440_ _0914_ _0917_ _0920_ VPWR VGND sg13g2_nor3_1
XFILLER_0_927 VPWR VGND sg13g2_decap_8
X_4319_ net684 VGND VPWR net231 u_usb_cdc.u_sie.in_byte_q\[2\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_28_666 VPWR VGND sg13g2_fill_2
XFILLER_42_124 VPWR VGND sg13g2_decap_4
XFILLER_15_338 VPWR VGND sg13g2_fill_1
XFILLER_23_360 VPWR VGND sg13g2_fill_1
XFILLER_3_710 VPWR VGND sg13g2_decap_8
XFILLER_3_787 VPWR VGND sg13g2_decap_8
Xfanout590 net592 net590 VPWR VGND sg13g2_buf_8
XFILLER_47_975 VPWR VGND sg13g2_decap_8
XFILLER_20_1015 VPWR VGND sg13g2_decap_8
XFILLER_34_603 VPWR VGND sg13g2_fill_1
X_3621_ VGND VPWR _0547_ _1511_ _1594_ _1917_ sg13g2_a21oi_1
X_3552_ _1528_ _0554_ _0560_ _0576_ VPWR VGND sg13g2_and3_2
X_2503_ net721 net757 _0739_ _0800_ VPWR VGND sg13g2_nor3_1
X_3483_ u_usb_cdc.u_sie.in_byte_q\[0\] u_usb_cdc.u_sie.in_byte_q\[1\] net230 _1477_
+ VPWR VGND sg13g2_a21o_1
X_2434_ _0732_ _0729_ _0731_ VPWR VGND sg13g2_nand2_1
X_2365_ _0548_ net783 net778 _0665_ VPWR VGND sg13g2_a21o_2
XFILLER_5_1009 VPWR VGND sg13g2_decap_8
X_4104_ net649 VGND VPWR net419 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[24\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2296_ net746 _0595_ _0598_ VPWR VGND sg13g2_nor2_1
XFILLER_38_942 VPWR VGND sg13g2_decap_8
X_4035_ net681 VGND VPWR net356 u_usb_cdc.u_sie.in_toggle_q\[2\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_24_113 VPWR VGND sg13g2_fill_1
XFILLER_40_639 VPWR VGND sg13g2_decap_8
XFILLER_21_831 VPWR VGND sg13g2_fill_1
XFILLER_21_853 VPWR VGND sg13g2_decap_4
X_3819_ _1750_ _1749_ net1007 VPWR VGND sg13g2_nand2b_1
XFILLER_21_897 VPWR VGND sg13g2_fill_1
XFILLER_4_507 VPWR VGND sg13g2_decap_8
XFILLER_0_724 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_decap_8
XFILLER_46_76 VPWR VGND sg13g2_fill_1
XFILLER_44_934 VPWR VGND sg13g2_decap_8
XFILLER_29_986 VPWR VGND sg13g2_decap_8
XFILLER_46_87 VPWR VGND sg13g2_fill_1
XFILLER_8_802 VPWR VGND sg13g2_fill_1
XFILLER_8_868 VPWR VGND sg13g2_decap_8
XFILLER_3_562 VPWR VGND sg13g2_decap_4
X_2150_ _0453_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] _1935_ VPWR VGND sg13g2_nand2_1
XFILLER_39_728 VPWR VGND sg13g2_decap_8
X_2081_ VPWR _1960_ u_usb_cdc.u_sie.u_phy_rx.state_q\[2\] VGND sg13g2_inv_1
XFILLER_47_772 VPWR VGND sg13g2_decap_8
XFILLER_34_444 VPWR VGND sg13g2_decap_4
XFILLER_35_978 VPWR VGND sg13g2_decap_8
XFILLER_15_691 VPWR VGND sg13g2_fill_2
XFILLER_34_499 VPWR VGND sg13g2_decap_4
X_2983_ _1132_ VPWR _0165_ VGND _1913_ _1130_ sg13g2_o21ai_1
X_3604_ _1577_ VPWR _1578_ VGND _1503_ _1571_ sg13g2_o21ai_1
X_3535_ _1511_ net716 net782 VPWR VGND sg13g2_nand2_1
X_3466_ net833 net832 net837 _1465_ VPWR VGND sg13g2_nor3_2
X_2417_ _0656_ net574 net715 _0715_ VPWR VGND sg13g2_nand3_1
X_3397_ net753 _1408_ _1419_ VPWR VGND sg13g2_nor2_1
XFILLER_29_216 VPWR VGND sg13g2_decap_8
X_2348_ VGND VPWR _0638_ net536 _0062_ _0648_ sg13g2_a21oi_1
X_2279_ net840 _1989_ _0581_ VPWR VGND sg13g2_and2_1
X_4018_ _0053_ net37 VPWR VGND sg13g2_buf_1
XFILLER_37_293 VPWR VGND sg13g2_decap_8
XFILLER_41_926 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_fill_2
XFILLER_12_149 VPWR VGND sg13g2_fill_2
XFILLER_21_650 VPWR VGND sg13g2_fill_1
XFILLER_5_827 VPWR VGND sg13g2_decap_8
XFILLER_0_521 VPWR VGND sg13g2_decap_8
XFILLER_0_598 VPWR VGND sg13g2_decap_8
XFILLER_48_569 VPWR VGND sg13g2_fill_2
XFILLER_48_558 VPWR VGND sg13g2_decap_8
XFILLER_17_901 VPWR VGND sg13g2_fill_1
XFILLER_31_403 VPWR VGND sg13g2_decap_8
XFILLER_31_447 VPWR VGND sg13g2_fill_1
XFILLER_40_970 VPWR VGND sg13g2_decap_8
Xhold109 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[14\] VPWR VGND
+ net151 sg13g2_dlygate4sd3_1
XFILLER_7_197 VPWR VGND sg13g2_fill_2
Xheichips25_usb_cdc_41 VPWR VGND uio_out[7] sg13g2_tielo
X_3320_ net335 net632 net1046 _1373_ VPWR VGND sg13g2_nand3_1
XFILLER_4_893 VPWR VGND sg13g2_decap_8
XFILLER_3_370 VPWR VGND sg13g2_decap_8
X_3251_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[28\] net816
+ _1319_ VPWR VGND sg13g2_nor2b_1
X_2202_ u_usb_cdc.u_sie.data_q\[3\] net548 _0504_ VPWR VGND sg13g2_xor2_1
X_3182_ VGND VPWR _1255_ _1257_ _1258_ net578 sg13g2_a21oi_1
XFILLER_39_503 VPWR VGND sg13g2_fill_2
X_2133_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\] u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\]
+ _2009_ VPWR VGND sg13g2_nor2b_1
X_2064_ VPWR _1943_ net444 VGND sg13g2_inv_1
X_2966_ _1049_ net825 _1054_ _1125_ VPWR VGND sg13g2_mux2_1
XFILLER_33_1014 VPWR VGND sg13g2_decap_8
X_2897_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net456 _1098_ _0113_ VPWR VGND sg13g2_mux2_1
Xhold610 _0164_ VPWR VGND net928 sg13g2_dlygate4sd3_1
Xhold621 u_usb_cdc.u_sie.phy_state_q\[4\] VPWR VGND net939 sg13g2_dlygate4sd3_1
Xhold632 _0010_ VPWR VGND net950 sg13g2_dlygate4sd3_1
Xhold654 _0005_ VPWR VGND net972 sg13g2_dlygate4sd3_1
Xhold643 _0254_ VPWR VGND net961 sg13g2_dlygate4sd3_1
Xhold676 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] VPWR VGND net994 sg13g2_dlygate4sd3_1
Xhold687 u_usb_cdc.u_sie.delay_cnt_q\[0\] VPWR VGND net1005 sg13g2_dlygate4sd3_1
Xhold665 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[2\] VPWR VGND
+ net983 sg13g2_dlygate4sd3_1
X_3518_ _1493_ VPWR _1494_ VGND net792 _1491_ sg13g2_o21ai_1
X_3449_ _1453_ net214 net580 VPWR VGND sg13g2_nand2_1
Xhold698 u_usb_cdc.sie_out_data\[3\] VPWR VGND net1016 sg13g2_dlygate4sd3_1
XFILLER_45_506 VPWR VGND sg13g2_fill_2
XFILLER_26_720 VPWR VGND sg13g2_decap_8
XFILLER_41_712 VPWR VGND sg13g2_decap_8
XFILLER_43_33 VPWR VGND sg13g2_fill_1
XFILLER_43_77 VPWR VGND sg13g2_fill_2
XFILLER_4_145 VPWR VGND sg13g2_fill_1
XFILLER_1_841 VPWR VGND sg13g2_decap_8
XFILLER_49_823 VPWR VGND sg13g2_decap_8
XFILLER_0_395 VPWR VGND sg13g2_decap_8
XFILLER_1_1023 VPWR VGND sg13g2_decap_4
XFILLER_16_230 VPWR VGND sg13g2_fill_2
XFILLER_16_285 VPWR VGND sg13g2_fill_1
XFILLER_20_907 VPWR VGND sg13g2_fill_2
X_2820_ net5 net1040 net637 _0078_ VPWR VGND sg13g2_mux2_1
XFILLER_31_266 VPWR VGND sg13g2_decap_8
XFILLER_31_277 VPWR VGND sg13g2_fill_2
XFILLER_9_952 VPWR VGND sg13g2_decap_8
XFILLER_13_992 VPWR VGND sg13g2_decap_8
X_2751_ VGND VPWR net833 _0528_ _0998_ _0997_ sg13g2_a21oi_1
X_2682_ _0948_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] _0947_ VPWR VGND sg13g2_nand2_1
X_4421_ net725 VGND VPWR net50 u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[0\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
X_4352_ net681 VGND VPWR _0354_ u_usb_cdc.sie_out_data\[7\] clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_4_690 VPWR VGND sg13g2_decap_8
X_4283_ net677 VGND VPWR _0285_ u_usb_cdc.u_ctrl_endp.rec_q\[1\] clknet_leaf_50_clk
+ sg13g2_dfrbpq_2
X_3303_ net301 net631 net1046 _1359_ VPWR VGND sg13g2_nand3_1
X_3234_ net805 net601 _1303_ _1304_ VPWR VGND sg13g2_nor3_1
X_3165_ _1240_ net814 _1241_ VPWR VGND sg13g2_xor2_1
X_3096_ _1203_ VPWR _0207_ VGND net708 _1151_ sg13g2_o21ai_1
X_2116_ _1992_ _1991_ net748 _1994_ VPWR VGND sg13g2_a21o_2
X_2047_ _1926_ net920 VPWR VGND sg13g2_inv_2
XFILLER_23_756 VPWR VGND sg13g2_decap_8
XFILLER_10_417 VPWR VGND sg13g2_fill_2
X_3998_ _1879_ net327 net316 VPWR VGND sg13g2_nand2_1
X_2949_ net483 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net603 _0144_ VPWR VGND sg13g2_mux2_1
Xhold451 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[59\] VPWR VGND
+ net493 sg13g2_dlygate4sd3_1
XFILLER_2_627 VPWR VGND sg13g2_decap_8
Xhold462 _0361_ VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold440 _0111_ VPWR VGND net482 sg13g2_dlygate4sd3_1
Xhold473 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[3\] VPWR VGND net515 sg13g2_dlygate4sd3_1
Xhold495 _0062_ VPWR VGND net537 sg13g2_dlygate4sd3_1
Xhold484 _0022_ VPWR VGND net526 sg13g2_dlygate4sd3_1
XFILLER_46_837 VPWR VGND sg13g2_decap_8
XFILLER_6_933 VPWR VGND sg13g2_decap_8
XFILLER_10_995 VPWR VGND sg13g2_decap_8
XFILLER_37_815 VPWR VGND sg13g2_fill_1
XFILLER_49_697 VPWR VGND sg13g2_decap_8
XFILLER_24_509 VPWR VGND sg13g2_fill_1
XFILLER_45_870 VPWR VGND sg13g2_decap_8
X_3921_ VGND VPWR net282 _1814_ _1815_ net622 sg13g2_a21oi_1
X_3852_ _1740_ _1772_ _1773_ _1774_ VPWR VGND sg13g2_nor3_1
X_2803_ net1066 net824 net828 _1044_ VPWR VGND u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ sg13g2_nand4_1
X_3783_ VPWR _0374_ net900 VGND sg13g2_inv_1
X_2734_ net745 _0595_ _0599_ _0981_ _0982_ VPWR VGND sg13g2_nor4_1
X_2665_ _0934_ _2012_ _0450_ VPWR VGND sg13g2_nand2_1
X_2596_ _0877_ u_usb_cdc.addr\[3\] net200 VPWR VGND sg13g2_xnor2_1
X_4404_ net728 VGND VPWR _0043_ u_usb_cdc.u_sie.u_phy_rx.rx_eop_q clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_4335_ net695 VGND VPWR net350 u_usb_cdc.u_sie.crc16_q\[14\] clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4266_ net679 VGND VPWR net270 u_usb_cdc.addr\[0\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_3217_ VGND VPWR _1274_ _1288_ _0243_ net405 sg13g2_a21oi_1
X_4197_ net661 VGND VPWR _0200_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[33\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3148_ _1231_ VPWR _0231_ VGND _1168_ _1229_ sg13g2_o21ai_1
X_3079_ _1194_ VPWR _0199_ VGND net721 net606 sg13g2_o21ai_1
XFILLER_35_380 VPWR VGND sg13g2_decap_4
XFILLER_24_35 VPWR VGND sg13g2_fill_1
XFILLER_10_214 VPWR VGND sg13g2_decap_8
XFILLER_10_247 VPWR VGND sg13g2_fill_1
XFILLER_7_719 VPWR VGND sg13g2_decap_8
XFILLER_2_413 VPWR VGND sg13g2_decap_8
Xhold270 _0059_ VPWR VGND net312 sg13g2_dlygate4sd3_1
XFILLER_6_4 VPWR VGND sg13g2_fill_2
XFILLER_3_969 VPWR VGND sg13g2_decap_8
XFILLER_49_32 VPWR VGND sg13g2_decap_8
Xhold281 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[52\] VPWR
+ VGND net323 sg13g2_dlygate4sd3_1
Xhold292 _0435_ VPWR VGND net334 sg13g2_dlygate4sd3_1
Xfanout750 net1044 net750 VPWR VGND sg13g2_buf_8
Xfanout761 net399 net761 VPWR VGND sg13g2_buf_8
Xfanout783 net784 net783 VPWR VGND sg13g2_buf_8
Xfanout772 net1031 net772 VPWR VGND sg13g2_buf_8
Xfanout794 net796 net794 VPWR VGND sg13g2_buf_8
XFILLER_45_122 VPWR VGND sg13g2_decap_8
XFILLER_46_689 VPWR VGND sg13g2_fill_1
XFILLER_41_383 VPWR VGND sg13g2_fill_1
XFILLER_14_586 VPWR VGND sg13g2_decap_4
XFILLER_6_730 VPWR VGND sg13g2_decap_8
X_2450_ VGND VPWR _0747_ u_usb_cdc.u_ctrl_endp.req_q\[11\] u_usb_cdc.u_ctrl_endp.req_q\[4\]
+ sg13g2_or2_1
X_2381_ _0605_ u_usb_cdc.u_ctrl_endp.state_q\[2\] _0681_ VPWR VGND sg13g2_nor2b_2
XFILLER_2_991 VPWR VGND sg13g2_decap_8
X_4120_ net655 VGND VPWR net84 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[40\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
X_4051_ net687 VGND VPWR _0026_ u_usb_cdc.u_sie.phy_state_q\[7\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_3002_ _1144_ net54 net614 VPWR VGND sg13g2_nand2_1
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
XFILLER_37_656 VPWR VGND sg13g2_decap_8
XFILLER_17_391 VPWR VGND sg13g2_decap_4
XFILLER_32_350 VPWR VGND sg13g2_decap_8
X_3904_ net929 net428 _0972_ _0416_ VPWR VGND sg13g2_mux2_1
XFILLER_33_851 VPWR VGND sg13g2_fill_2
XFILLER_33_873 VPWR VGND sg13g2_decap_8
XFILLER_20_501 VPWR VGND sg13g2_fill_2
XFILLER_32_383 VPWR VGND sg13g2_fill_2
X_3835_ _1761_ net710 net402 VPWR VGND sg13g2_nand2_1
XFILLER_20_556 VPWR VGND sg13g2_fill_1
X_3766_ _1710_ VPWR _1711_ VGND net833 _1709_ sg13g2_o21ai_1
X_2717_ net703 _0939_ _0972_ VPWR VGND sg13g2_nor2_2
X_3697_ _1666_ net491 _1360_ VPWR VGND sg13g2_nand2_1
X_2648_ _0919_ _0441_ _0917_ VPWR VGND sg13g2_nand2_1
XFILLER_0_906 VPWR VGND sg13g2_decap_8
X_2579_ VPWR VGND _0862_ _0646_ _0856_ _0554_ _0863_ _0638_ sg13g2_a221oi_1
X_4318_ net683 VGND VPWR net320 u_usb_cdc.u_sie.in_byte_q\[1\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_4249_ net653 VGND VPWR net969 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[1\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_2
XFILLER_28_634 VPWR VGND sg13g2_decap_4
XFILLER_43_604 VPWR VGND sg13g2_fill_2
XFILLER_35_67 VPWR VGND sg13g2_fill_1
XFILLER_11_578 VPWR VGND sg13g2_fill_1
XFILLER_3_766 VPWR VGND sg13g2_decap_8
XFILLER_2_287 VPWR VGND sg13g2_fill_2
Xfanout580 net582 net580 VPWR VGND sg13g2_buf_8
Xfanout591 net592 net591 VPWR VGND sg13g2_buf_1
XFILLER_47_954 VPWR VGND sg13g2_decap_8
XFILLER_19_656 VPWR VGND sg13g2_decap_8
XFILLER_15_851 VPWR VGND sg13g2_fill_1
XFILLER_30_854 VPWR VGND sg13g2_fill_1
X_3620_ net773 _0669_ _1593_ VPWR VGND sg13g2_nor2_1
X_3551_ _1523_ _1526_ _1522_ _1527_ VPWR VGND sg13g2_nand3_1
X_2502_ VPWR _0799_ _0798_ VGND sg13g2_inv_1
X_3482_ _1476_ net230 net594 VPWR VGND sg13g2_nand2_1
X_2433_ net760 net757 _0730_ _0731_ VPWR VGND sg13g2_nor3_1
X_2364_ _0664_ net786 net780 VPWR VGND sg13g2_nand2_1
X_4103_ net668 VGND VPWR net68 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[23\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_2295_ _0597_ net208 net595 VPWR VGND sg13g2_nand2_1
XFILLER_38_921 VPWR VGND sg13g2_decap_8
X_4034_ net681 VGND VPWR net925 u_usb_cdc.u_sie.in_toggle_q\[1\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_37_464 VPWR VGND sg13g2_decap_8
XFILLER_38_998 VPWR VGND sg13g2_decap_8
XFILLER_24_103 VPWR VGND sg13g2_fill_1
XFILLER_24_169 VPWR VGND sg13g2_fill_2
XFILLER_40_607 VPWR VGND sg13g2_decap_4
XFILLER_21_821 VPWR VGND sg13g2_fill_2
XFILLER_32_191 VPWR VGND sg13g2_decap_4
X_3818_ net318 net331 net740 _1749_ VPWR VGND net202 sg13g2_nand4_1
X_3749_ net904 _1697_ _1695_ _0366_ VPWR VGND sg13g2_mux2_1
XFILLER_0_703 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_43_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_228 VPWR VGND sg13g2_decap_4
XFILLER_29_965 VPWR VGND sg13g2_decap_8
XFILLER_44_913 VPWR VGND sg13g2_decap_8
XFILLER_43_456 VPWR VGND sg13g2_fill_1
XFILLER_43_445 VPWR VGND sg13g2_fill_2
XFILLER_24_670 VPWR VGND sg13g2_decap_8
XFILLER_11_320 VPWR VGND sg13g2_decap_8
XFILLER_12_887 VPWR VGND sg13g2_fill_1
XFILLER_3_552 VPWR VGND sg13g2_fill_1
XFILLER_38_206 VPWR VGND sg13g2_decap_8
XFILLER_47_751 VPWR VGND sg13g2_decap_8
X_2080_ VPWR _1959_ net189 VGND sg13g2_inv_1
XFILLER_19_475 VPWR VGND sg13g2_decap_8
XFILLER_19_486 VPWR VGND sg13g2_fill_1
XFILLER_19_497 VPWR VGND sg13g2_fill_2
XFILLER_34_423 VPWR VGND sg13g2_decap_8
XFILLER_35_957 VPWR VGND sg13g2_decap_8
XFILLER_34_456 VPWR VGND sg13g2_decap_8
X_2982_ _1132_ net280 _1130_ VPWR VGND sg13g2_nand2_1
XFILLER_21_106 VPWR VGND sg13g2_fill_1
XFILLER_30_662 VPWR VGND sg13g2_fill_1
X_3603_ VGND VPWR net770 _1576_ _1577_ _1516_ sg13g2_a21oi_1
X_3534_ net777 _0547_ _1510_ VPWR VGND sg13g2_and2_1
X_3465_ _1464_ _0494_ _1463_ _0315_ VPWR VGND sg13g2_a21o_1
X_2416_ _0714_ net760 _0709_ VPWR VGND sg13g2_nand2_1
X_3396_ net854 net567 _1418_ VPWR VGND sg13g2_nor2_1
X_2347_ _0645_ VPWR _0648_ VGND net535 _0647_ sg13g2_o21ai_1
X_2278_ _0580_ net839 _0579_ VPWR VGND sg13g2_nand2_1
XFILLER_38_762 VPWR VGND sg13g2_fill_2
XFILLER_38_784 VPWR VGND sg13g2_decap_4
X_4017_ VPWR _0439_ net565 VGND sg13g2_inv_1
XFILLER_41_905 VPWR VGND sg13g2_decap_8
XFILLER_25_456 VPWR VGND sg13g2_decap_8
XFILLER_12_106 VPWR VGND sg13g2_fill_2
XFILLER_13_618 VPWR VGND sg13g2_decap_4
XFILLER_5_806 VPWR VGND sg13g2_decap_8
XFILLER_0_500 VPWR VGND sg13g2_decap_8
XFILLER_0_577 VPWR VGND sg13g2_decap_8
XFILLER_48_537 VPWR VGND sg13g2_decap_8
XFILLER_44_732 VPWR VGND sg13g2_fill_2
XFILLER_16_401 VPWR VGND sg13g2_fill_1
XFILLER_16_412 VPWR VGND sg13g2_decap_8
XFILLER_16_423 VPWR VGND sg13g2_fill_2
XFILLER_28_294 VPWR VGND sg13g2_decap_8
XFILLER_44_798 VPWR VGND sg13g2_decap_4
XFILLER_12_651 VPWR VGND sg13g2_fill_1
XFILLER_8_688 VPWR VGND sg13g2_fill_1
XFILLER_7_187 VPWR VGND sg13g2_fill_2
XFILLER_4_872 VPWR VGND sg13g2_decap_8
X_3250_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[4\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[12\]
+ net816 _1318_ VPWR VGND sg13g2_mux2_1
XFILLER_26_1022 VPWR VGND sg13g2_decap_8
X_2201_ _0503_ _0501_ _0502_ VPWR VGND sg13g2_xnor2_1
X_3181_ _1257_ _0606_ _1256_ net955 net749 VPWR VGND sg13g2_a22oi_1
X_2132_ net988 net973 _2008_ VPWR VGND sg13g2_nor2b_2
XFILLER_39_548 VPWR VGND sg13g2_fill_1
X_2063_ VPWR _1942_ u_usb_cdc.u_sie.crc16_q\[11\] VGND sg13g2_inv_1
XFILLER_23_949 VPWR VGND sg13g2_fill_1
XFILLER_34_253 VPWR VGND sg13g2_fill_1
XFILLER_22_437 VPWR VGND sg13g2_decap_8
X_2965_ net870 _1124_ _1123_ _0155_ VPWR VGND sg13g2_mux2_1
XFILLER_31_982 VPWR VGND sg13g2_decap_8
X_2896_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net410 _1098_ _0112_ VPWR VGND sg13g2_mux2_1
Xhold600 u_usb_cdc.u_sie.crc16_q\[1\] VPWR VGND net918 sg13g2_dlygate4sd3_1
Xhold611 u_usb_cdc.u_sie.rx_data\[4\] VPWR VGND net929 sg13g2_dlygate4sd3_1
XFILLER_2_809 VPWR VGND sg13g2_decap_8
Xhold633 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] VPWR VGND net951 sg13g2_dlygate4sd3_1
Xhold622 u_usb_cdc.u_sie.rx_data\[1\] VPWR VGND net940 sg13g2_dlygate4sd3_1
Xhold644 net27 VPWR VGND net962 sg13g2_dlygate4sd3_1
X_3517_ VGND VPWR net792 _1492_ _1493_ net789 sg13g2_a21oi_1
Xhold655 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[0\] VPWR VGND net973 sg13g2_dlygate4sd3_1
Xhold688 _0316_ VPWR VGND net1006 sg13g2_dlygate4sd3_1
Xhold666 _0253_ VPWR VGND net984 sg13g2_dlygate4sd3_1
Xhold677 u_usb_cdc.u_sie.data_q\[5\] VPWR VGND net995 sg13g2_dlygate4sd3_1
X_3448_ _1452_ VPWR _0310_ VGND _1899_ net581 sg13g2_o21ai_1
Xhold699 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\] VPWR
+ VGND net1017 sg13g2_dlygate4sd3_1
X_3379_ _0724_ _1405_ _1406_ VPWR VGND sg13g2_nor2_1
XFILLER_40_1019 VPWR VGND sg13g2_decap_8
XFILLER_25_220 VPWR VGND sg13g2_decap_4
XFILLER_26_776 VPWR VGND sg13g2_fill_1
XFILLER_9_408 VPWR VGND sg13g2_fill_2
XFILLER_13_426 VPWR VGND sg13g2_decap_8
XFILLER_13_448 VPWR VGND sg13g2_decap_4
XFILLER_43_89 VPWR VGND sg13g2_fill_1
XFILLER_5_647 VPWR VGND sg13g2_fill_1
XFILLER_1_820 VPWR VGND sg13g2_decap_8
XFILLER_49_802 VPWR VGND sg13g2_decap_8
XFILLER_1_897 VPWR VGND sg13g2_decap_8
XFILLER_0_374 VPWR VGND sg13g2_decap_8
XFILLER_49_879 VPWR VGND sg13g2_decap_8
XFILLER_1_1002 VPWR VGND sg13g2_decap_8
XFILLER_17_90 VPWR VGND sg13g2_fill_1
XFILLER_13_971 VPWR VGND sg13g2_decap_8
XFILLER_8_430 VPWR VGND sg13g2_fill_1
XFILLER_9_931 VPWR VGND sg13g2_decap_8
X_2750_ _0604_ _0996_ _0590_ _0997_ VPWR VGND sg13g2_nand3_1
XFILLER_8_452 VPWR VGND sg13g2_fill_1
X_2681_ net711 _1959_ _0947_ VPWR VGND sg13g2_nor2_1
X_4420_ net729 VGND VPWR net361 u_usb_cdc.u_sie.rx_data\[7\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_4351_ net681 VGND VPWR _0353_ u_usb_cdc.sie_out_data\[6\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_4282_ net665 VGND VPWR _0284_ u_usb_cdc.u_ctrl_endp.rec_q\[0\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_2
X_3302_ _1358_ _1123_ _1129_ VPWR VGND sg13g2_nand2_2
X_3233_ VPWR VGND _1279_ _1301_ _1302_ net808 _1303_ _1298_ sg13g2_a221oi_1
XFILLER_39_334 VPWR VGND sg13g2_fill_2
X_3164_ VGND VPWR net1070 _1148_ _1240_ net822 sg13g2_a21oi_1
X_3095_ _1203_ net78 _1202_ VPWR VGND sg13g2_nand2_1
XFILLER_27_529 VPWR VGND sg13g2_fill_2
X_2115_ VGND VPWR net747 _1993_ _1992_ _1991_ sg13g2_a21oi_2
XFILLER_35_540 VPWR VGND sg13g2_fill_1
X_2046_ _1925_ u_usb_cdc.u_sie.pid_q\[3\] VPWR VGND sg13g2_inv_2
X_3997_ _1878_ net316 net713 VPWR VGND sg13g2_nand2_1
X_2948_ net487 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ _1119_ _0143_ VPWR VGND sg13g2_mux2_1
X_2879_ _1091_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ _1082_ VPWR VGND sg13g2_nand2_1
XFILLER_2_606 VPWR VGND sg13g2_decap_8
Xhold441 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[61\] VPWR VGND
+ net483 sg13g2_dlygate4sd3_1
Xhold452 _0142_ VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold463 net17 VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold430 _0116_ VPWR VGND net472 sg13g2_dlygate4sd3_1
Xhold496 u_usb_cdc.u_ctrl_endp.max_length_q\[4\] VPWR VGND net538 sg13g2_dlygate4sd3_1
Xhold474 _1735_ VPWR VGND net516 sg13g2_dlygate4sd3_1
Xhold485 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[4\] VPWR VGND net527 sg13g2_dlygate4sd3_1
XFILLER_46_816 VPWR VGND sg13g2_decap_8
XFILLER_13_223 VPWR VGND sg13g2_decap_8
XFILLER_41_598 VPWR VGND sg13g2_fill_2
XFILLER_6_912 VPWR VGND sg13g2_decap_8
XFILLER_10_974 VPWR VGND sg13g2_decap_8
XFILLER_6_989 VPWR VGND sg13g2_decap_8
XFILLER_49_632 VPWR VGND sg13g2_decap_4
XFILLER_1_694 VPWR VGND sg13g2_decap_8
XFILLER_49_676 VPWR VGND sg13g2_decap_8
XFILLER_17_551 VPWR VGND sg13g2_decap_8
XFILLER_17_562 VPWR VGND sg13g2_fill_1
X_3920_ _1994_ _1034_ _1814_ VPWR VGND sg13g2_nor2_1
XFILLER_44_381 VPWR VGND sg13g2_decap_4
X_3851_ _1773_ net422 net887 _1768_ VPWR VGND sg13g2_and3_1
X_2802_ _1043_ net828 net827 VPWR VGND sg13g2_nand2_2
X_3782_ _1723_ _1720_ net899 net579 net485 VPWR VGND sg13g2_a22oi_1
X_2733_ u_usb_cdc.u_sie.phy_state_q\[8\] net832 _0981_ VPWR VGND sg13g2_nor2_1
X_2664_ _0932_ net935 net703 _0933_ VPWR VGND sg13g2_a21o_2
X_2595_ u_usb_cdc.u_sie.addr_q\[5\] u_usb_cdc.addr\[5\] _0876_ VPWR VGND sg13g2_xor2_1
X_4403_ net725 VGND VPWR net936 u_usb_cdc.u_sie.u_phy_rx.rx_en_q clknet_leaf_39_clk
+ sg13g2_dfrbpq_2
X_4334_ net687 VGND VPWR net307 u_usb_cdc.u_sie.crc16_q\[13\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_8_1008 VPWR VGND sg13g2_decap_8
X_4265_ net676 VGND VPWR net480 u_usb_cdc.u_ctrl_endp.in_endp_q clknet_leaf_44_clk
+ sg13g2_dfrbpq_2
X_3216_ VGND VPWR net118 _1287_ _1288_ _1285_ sg13g2_a21oi_1
X_4196_ net665 VGND VPWR net243 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[32\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3147_ _1231_ net118 _1230_ VPWR VGND sg13g2_nand2_1
XFILLER_27_304 VPWR VGND sg13g2_fill_1
XFILLER_27_359 VPWR VGND sg13g2_fill_2
X_3078_ _1194_ net242 net606 VPWR VGND sg13g2_nand2_1
X_2029_ VPWR _1908_ net964 VGND sg13g2_inv_1
XFILLER_23_510 VPWR VGND sg13g2_fill_2
XFILLER_10_204 VPWR VGND sg13g2_fill_1
XFILLER_6_219 VPWR VGND sg13g2_fill_2
XFILLER_49_11 VPWR VGND sg13g2_decap_8
Xhold260 _0163_ VPWR VGND net302 sg13g2_dlygate4sd3_1
Xhold271 _0430_ VPWR VGND net313 sg13g2_dlygate4sd3_1
XFILLER_3_948 VPWR VGND sg13g2_decap_8
Xhold282 _0219_ VPWR VGND net324 sg13g2_dlygate4sd3_1
XFILLER_2_469 VPWR VGND sg13g2_decap_8
Xhold293 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[3\] VPWR VGND
+ net335 sg13g2_dlygate4sd3_1
Xfanout740 net742 net740 VPWR VGND sg13g2_buf_8
Xfanout751 net942 net751 VPWR VGND sg13g2_buf_8
Xfanout784 net1060 net784 VPWR VGND sg13g2_buf_8
Xfanout773 net775 net773 VPWR VGND sg13g2_buf_8
Xfanout762 net763 net762 VPWR VGND sg13g2_buf_8
Xfanout795 net796 net795 VPWR VGND sg13g2_buf_1
XFILLER_46_657 VPWR VGND sg13g2_fill_1
XFILLER_27_860 VPWR VGND sg13g2_fill_1
XFILLER_6_786 VPWR VGND sg13g2_decap_8
XFILLER_2_970 VPWR VGND sg13g2_decap_8
X_2380_ VGND VPWR _0680_ net588 net714 sg13g2_or2_1
XFILLER_39_5 VPWR VGND sg13g2_decap_8
XFILLER_1_491 VPWR VGND sg13g2_decap_8
X_4050_ net697 VGND VPWR net209 u_usb_cdc.u_sie.phy_state_q\[6\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
XFILLER_49_484 VPWR VGND sg13g2_decap_8
X_3001_ _1143_ VPWR _0172_ VGND _1898_ net613 sg13g2_o21ai_1
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
XFILLER_37_624 VPWR VGND sg13g2_fill_1
XFILLER_17_370 VPWR VGND sg13g2_fill_1
XFILLER_33_830 VPWR VGND sg13g2_decap_8
X_3903_ net966 net527 net599 _0415_ VPWR VGND sg13g2_mux2_1
X_3834_ net873 net710 _1760_ _0388_ VPWR VGND sg13g2_a21o_1
XFILLER_32_395 VPWR VGND sg13g2_fill_2
X_3765_ VGND VPWR _1466_ _1709_ _1710_ net712 sg13g2_a21oi_1
X_2716_ VGND VPWR net704 _0971_ _0047_ _0970_ sg13g2_a21oi_1
X_3696_ _1665_ net919 net593 VPWR VGND sg13g2_nand2_1
X_2647_ _0914_ VPWR _0918_ VGND u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\] u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[0\]
+ sg13g2_o21ai_1
X_2578_ u_usb_cdc.sie_in_data_ack _0554_ net583 _0862_ VPWR VGND sg13g2_nor3_1
X_4317_ net684 VGND VPWR net290 u_usb_cdc.u_sie.in_byte_q\[0\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
X_4248_ net653 VGND VPWR net956 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[0\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_2
XFILLER_28_624 VPWR VGND sg13g2_decap_4
X_4179_ net646 VGND VPWR net222 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[15\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_43_638 VPWR VGND sg13g2_decap_4
XFILLER_15_329 VPWR VGND sg13g2_decap_8
XFILLER_23_373 VPWR VGND sg13g2_decap_8
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_13_1013 VPWR VGND sg13g2_decap_8
XFILLER_3_745 VPWR VGND sg13g2_decap_8
XFILLER_2_222 VPWR VGND sg13g2_fill_2
XFILLER_47_933 VPWR VGND sg13g2_decap_8
Xfanout570 _1388_ net570 VPWR VGND sg13g2_buf_8
Xfanout581 net582 net581 VPWR VGND sg13g2_buf_1
XFILLER_19_602 VPWR VGND sg13g2_fill_2
Xfanout592 _0594_ net592 VPWR VGND sg13g2_buf_8
XFILLER_14_362 VPWR VGND sg13g2_fill_1
XFILLER_30_800 VPWR VGND sg13g2_fill_2
X_3550_ _1526_ _1525_ _1524_ VPWR VGND sg13g2_nand2b_1
X_2501_ net920 net910 net993 _0798_ VPWR VGND sg13g2_nor3_1
X_3481_ _1474_ VPWR _0320_ VGND _0894_ _1475_ sg13g2_o21ai_1
X_2432_ net718 _0707_ net1016 _0730_ VPWR VGND sg13g2_nand3_1
X_2363_ _0656_ _0659_ net715 _0663_ VPWR VGND sg13g2_nand3_1
X_4102_ net669 VGND VPWR net148 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[22\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
X_4033_ net691 VGND VPWR net311 u_usb_cdc.u_sie.in_toggle_q\[0\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_2294_ net260 net592 _0580_ _0596_ VPWR VGND sg13g2_nand3_1
XFILLER_38_911 VPWR VGND sg13g2_fill_1
XFILLER_37_443 VPWR VGND sg13g2_decap_8
XFILLER_38_977 VPWR VGND sg13g2_decap_8
XFILLER_18_690 VPWR VGND sg13g2_fill_2
XFILLER_36_1024 VPWR VGND sg13g2_decap_4
X_3817_ net740 VPWR _1748_ VGND _1738_ _1747_ sg13g2_o21ai_1
XFILLER_21_888 VPWR VGND sg13g2_decap_8
X_3748_ _1696_ VPWR _1697_ VGND _0890_ _1693_ sg13g2_o21ai_1
X_3679_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[22\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[30\]
+ net800 _1649_ VPWR VGND sg13g2_mux2_1
XFILLER_43_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_759 VPWR VGND sg13g2_decap_8
XFILLER_28_410 VPWR VGND sg13g2_decap_8
XFILLER_15_115 VPWR VGND sg13g2_fill_2
XFILLER_16_638 VPWR VGND sg13g2_fill_2
XFILLER_44_969 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_50_clk clknet_3_1__leaf_clk clknet_leaf_50_clk VPWR VGND sg13g2_buf_8
XFILLER_8_826 VPWR VGND sg13g2_fill_2
XFILLER_11_398 VPWR VGND sg13g2_fill_1
XFILLER_3_597 VPWR VGND sg13g2_fill_2
XFILLER_3_586 VPWR VGND sg13g2_decap_8
XFILLER_23_8 VPWR VGND sg13g2_decap_4
XFILLER_47_730 VPWR VGND sg13g2_decap_8
XFILLER_19_465 VPWR VGND sg13g2_fill_1
XFILLER_35_936 VPWR VGND sg13g2_decap_8
X_2981_ net794 net927 _1130_ _0164_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_41_clk clknet_3_5__leaf_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
XFILLER_30_652 VPWR VGND sg13g2_fill_2
X_3602_ VGND VPWR _0650_ _1429_ _1576_ _1575_ sg13g2_a21oi_1
XFILLER_30_685 VPWR VGND sg13g2_decap_4
XFILLER_7_892 VPWR VGND sg13g2_decap_8
X_3533_ _1502_ VPWR _1509_ VGND _1506_ _1508_ sg13g2_o21ai_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_3464_ _0589_ _0591_ _0976_ _1464_ VPWR VGND sg13g2_nor3_1
X_2415_ net721 _0710_ _0713_ VPWR VGND sg13g2_nor2_2
X_3395_ VGND VPWR net568 _1417_ _0292_ _1416_ sg13g2_a21oi_1
X_2346_ _0647_ _0646_ VPWR VGND sg13g2_inv_2
X_2277_ _0579_ _0578_ VPWR VGND _0577_ sg13g2_nand2b_2
X_4016_ _1891_ VPWR _1892_ VGND net737 net564 sg13g2_o21ai_1
XFILLER_38_752 VPWR VGND sg13g2_fill_1
XFILLER_25_402 VPWR VGND sg13g2_decap_8
XFILLER_16_48 VPWR VGND sg13g2_decap_4
XFILLER_34_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_32_clk clknet_3_7__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_20_140 VPWR VGND sg13g2_decap_4
XFILLER_21_696 VPWR VGND sg13g2_fill_2
XFILLER_10_1016 VPWR VGND sg13g2_decap_8
XFILLER_10_1027 VPWR VGND sg13g2_fill_2
XFILLER_0_556 VPWR VGND sg13g2_decap_8
XFILLER_48_516 VPWR VGND sg13g2_decap_8
XFILLER_44_722 VPWR VGND sg13g2_fill_1
XFILLER_28_262 VPWR VGND sg13g2_fill_2
XFILLER_28_273 VPWR VGND sg13g2_decap_8
XFILLER_44_744 VPWR VGND sg13g2_fill_2
XFILLER_16_435 VPWR VGND sg13g2_decap_8
XFILLER_16_468 VPWR VGND sg13g2_decap_8
XFILLER_43_298 VPWR VGND sg13g2_fill_2
XFILLER_24_490 VPWR VGND sg13g2_fill_2
XFILLER_31_438 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_23_clk clknet_3_6__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_4_851 VPWR VGND sg13g2_decap_8
X_2200_ u_usb_cdc.u_sie.data_q\[5\] net444 _0502_ VPWR VGND sg13g2_xor2_1
XFILLER_26_1001 VPWR VGND sg13g2_decap_8
X_3180_ net822 net955 net768 _1256_ VPWR VGND sg13g2_mux2_1
XFILLER_39_505 VPWR VGND sg13g2_fill_1
X_2131_ _0065_ net712 _1983_ VPWR VGND sg13g2_nand2_1
X_2062_ VPWR _1941_ u_usb_cdc.u_sie.crc16_q\[12\] VGND sg13g2_inv_1
XFILLER_34_221 VPWR VGND sg13g2_decap_4
XFILLER_22_416 VPWR VGND sg13g2_decap_8
X_2964_ _1045_ net827 _1054_ _1124_ VPWR VGND sg13g2_mux2_1
XFILLER_34_298 VPWR VGND sg13g2_fill_2
XFILLER_31_961 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_14_clk clknet_3_2__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_2895_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net481 _1098_ _0111_ VPWR VGND sg13g2_mux2_1
Xhold612 _0416_ VPWR VGND net930 sg13g2_dlygate4sd3_1
Xhold601 u_usb_cdc.u_sie.data_q\[7\] VPWR VGND net919 sg13g2_dlygate4sd3_1
Xhold634 _0301_ VPWR VGND net952 sg13g2_dlygate4sd3_1
Xhold645 _0364_ VPWR VGND net963 sg13g2_dlygate4sd3_1
Xhold623 u_usb_cdc.in_ready_o[0] VPWR VGND net941 sg13g2_dlygate4sd3_1
X_3516_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[16\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[24\]
+ net797 _1492_ VPWR VGND sg13g2_mux2_1
Xhold678 u_usb_cdc.sie_out_data\[4\] VPWR VGND net996 sg13g2_dlygate4sd3_1
Xhold656 _0407_ VPWR VGND net974 sg13g2_dlygate4sd3_1
Xhold667 u_usb_cdc.u_sie.data_q\[6\] VPWR VGND net985 sg13g2_dlygate4sd3_1
Xhold689 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[3\] VPWR VGND net1007 sg13g2_dlygate4sd3_1
X_3447_ _1452_ net237 net581 VPWR VGND sg13g2_nand2_1
X_3378_ net620 _0675_ _1404_ _1405_ VPWR VGND sg13g2_nor3_1
X_2329_ VGND VPWR _1909_ net841 _0630_ u_usb_cdc.u_ctrl_endp.state_q\[2\] sg13g2_a21oi_1
XFILLER_45_508 VPWR VGND sg13g2_fill_1
XFILLER_27_58 VPWR VGND sg13g2_decap_8
XFILLER_13_416 VPWR VGND sg13g2_fill_1
XFILLER_43_79 VPWR VGND sg13g2_fill_1
XFILLER_21_460 VPWR VGND sg13g2_fill_2
XFILLER_21_471 VPWR VGND sg13g2_fill_1
XFILLER_49_1012 VPWR VGND sg13g2_decap_8
XFILLER_4_136 VPWR VGND sg13g2_decap_8
XFILLER_0_353 VPWR VGND sg13g2_decap_8
XFILLER_1_876 VPWR VGND sg13g2_decap_8
XFILLER_49_858 VPWR VGND sg13g2_decap_8
XFILLER_17_788 VPWR VGND sg13g2_fill_1
XFILLER_31_202 VPWR VGND sg13g2_fill_2
XFILLER_9_910 VPWR VGND sg13g2_decap_8
XFILLER_13_950 VPWR VGND sg13g2_decap_8
XFILLER_20_909 VPWR VGND sg13g2_fill_1
XFILLER_12_460 VPWR VGND sg13g2_fill_1
XFILLER_9_987 VPWR VGND sg13g2_decap_8
X_2680_ _0945_ VPWR _0032_ VGND _0913_ _0946_ sg13g2_o21ai_1
XFILLER_8_486 VPWR VGND sg13g2_decap_8
X_4350_ net691 VGND VPWR _0352_ u_usb_cdc.sie_out_data\[5\] clknet_leaf_46_clk sg13g2_dfrbpq_2
X_3301_ _1296_ _1357_ _0258_ VPWR VGND sg13g2_nor2_1
X_4281_ net679 VGND VPWR _0283_ u_usb_cdc.u_ctrl_endp.dev_state_q\[1\] clknet_leaf_47_clk
+ sg13g2_dfrbpq_1
X_3232_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[2\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[10\]
+ net817 _1302_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3163_ net633 _0609_ net739 _1239_ VPWR VGND sg13g2_nand3_1
XFILLER_39_324 VPWR VGND sg13g2_fill_1
X_2114_ net838 net834 u_usb_cdc.u_sie.phy_state_q\[11\] net831 _1992_ VPWR VGND sg13g2_nor4_1
XFILLER_39_346 VPWR VGND sg13g2_decap_8
XFILLER_39_368 VPWR VGND sg13g2_fill_2
X_3094_ net822 net820 net737 _1202_ VPWR VGND _1134_ sg13g2_nand4_1
XFILLER_27_519 VPWR VGND sg13g2_fill_1
X_2045_ _1924_ u_usb_cdc.u_sie.pid_q\[2\] VPWR VGND sg13g2_inv_2
XFILLER_22_268 VPWR VGND sg13g2_decap_8
X_3996_ _1877_ VPWR _0433_ VGND net327 _1876_ sg13g2_o21ai_1
X_2947_ net493 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net603 _0142_ VPWR VGND sg13g2_mux2_1
XFILLER_10_419 VPWR VGND sg13g2_fill_1
XFILLER_13_38 VPWR VGND sg13g2_fill_2
X_2878_ _1090_ net61 _1080_ VPWR VGND sg13g2_nand2_1
Xhold420 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[62\] VPWR VGND
+ net462 sg13g2_dlygate4sd3_1
Xhold442 _0144_ VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold453 net31 VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold431 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[31\] VPWR VGND
+ net473 sg13g2_dlygate4sd3_1
Xhold464 _0358_ VPWR VGND net506 sg13g2_dlygate4sd3_1
Xhold486 _1724_ VPWR VGND net528 sg13g2_dlygate4sd3_1
Xhold475 _0380_ VPWR VGND net517 sg13g2_dlygate4sd3_1
Xhold497 _0292_ VPWR VGND net539 sg13g2_dlygate4sd3_1
XFILLER_14_769 VPWR VGND sg13g2_decap_4
XFILLER_10_953 VPWR VGND sg13g2_decap_8
XFILLER_6_968 VPWR VGND sg13g2_decap_8
XFILLER_1_673 VPWR VGND sg13g2_decap_8
XFILLER_23_1004 VPWR VGND sg13g2_decap_4
XFILLER_49_655 VPWR VGND sg13g2_decap_8
XFILLER_23_1026 VPWR VGND sg13g2_fill_2
XFILLER_36_327 VPWR VGND sg13g2_fill_2
XFILLER_17_541 VPWR VGND sg13g2_fill_1
XFILLER_32_511 VPWR VGND sg13g2_decap_8
XFILLER_32_522 VPWR VGND sg13g2_fill_2
X_3850_ VGND VPWR net422 _1768_ _1772_ net887 sg13g2_a21oi_1
XFILLER_32_555 VPWR VGND sg13g2_fill_2
X_2801_ _1042_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[0\] _1041_
+ VPWR VGND sg13g2_xnor2_1
X_3781_ VPWR _0373_ net486 VGND sg13g2_inv_1
XFILLER_32_577 VPWR VGND sg13g2_fill_2
XFILLER_13_791 VPWR VGND sg13g2_decap_8
X_2732_ _0980_ _0979_ _0494_ _0601_ _0498_ VPWR VGND sg13g2_a22oi_1
XFILLER_8_250 VPWR VGND sg13g2_fill_1
XFILLER_30_1019 VPWR VGND sg13g2_decap_4
XFILLER_8_283 VPWR VGND sg13g2_fill_2
X_2663_ _0930_ _0931_ _0932_ VPWR VGND sg13g2_nor2_1
X_2594_ _0875_ u_usb_cdc.addr\[1\] net252 VPWR VGND sg13g2_xnor2_1
X_4402_ net728 VGND VPWR _0404_ u_usb_cdc.u_sie.rx_err clknet_leaf_33_clk sg13g2_dfrbpq_1
X_4333_ net687 VGND VPWR net286 u_usb_cdc.u_sie.crc16_q\[12\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_5_72 VPWR VGND sg13g2_decap_8
X_4264_ net676 VGND VPWR _0266_ u_usb_cdc.u_ctrl_endp.endp_q\[3\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
X_3215_ net812 _1286_ _1287_ VPWR VGND sg13g2_nor2_1
X_4195_ net662 VGND VPWR _0198_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[31\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3146_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\] _1148_
+ net735 _1230_ VPWR VGND sg13g2_nand3_1
X_3077_ _1134_ _1136_ net820 _1193_ VPWR VGND sg13g2_nand3_1
XFILLER_42_319 VPWR VGND sg13g2_decap_8
X_2028_ VPWR _1907_ net958 VGND sg13g2_inv_1
XFILLER_23_533 VPWR VGND sg13g2_fill_2
XFILLER_39_1022 VPWR VGND sg13g2_decap_8
XFILLER_35_393 VPWR VGND sg13g2_fill_2
X_3979_ _1863_ _1864_ _1993_ _1866_ VPWR VGND _1865_ sg13g2_nand4_1
XFILLER_3_927 VPWR VGND sg13g2_decap_8
XFILLER_2_448 VPWR VGND sg13g2_decap_8
Xhold261 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[10\] VPWR VGND net303 sg13g2_dlygate4sd3_1
Xhold250 _1717_ VPWR VGND net292 sg13g2_dlygate4sd3_1
XFILLER_46_1026 VPWR VGND sg13g2_fill_2
Xhold283 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[51\] VPWR
+ VGND net325 sg13g2_dlygate4sd3_1
Xhold272 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[23\] VPWR
+ VGND net314 sg13g2_dlygate4sd3_1
Xhold294 _0166_ VPWR VGND net336 sg13g2_dlygate4sd3_1
Xfanout741 net742 net741 VPWR VGND sg13g2_buf_8
Xfanout730 net731 net730 VPWR VGND sg13g2_buf_8
Xfanout752 net991 net752 VPWR VGND sg13g2_buf_8
Xfanout785 net1043 net785 VPWR VGND sg13g2_buf_8
Xfanout774 net775 net774 VPWR VGND sg13g2_buf_1
Xfanout763 net1023 net763 VPWR VGND sg13g2_buf_8
Xfanout796 net1026 net796 VPWR VGND sg13g2_buf_8
XFILLER_42_875 VPWR VGND sg13g2_fill_2
XFILLER_42_886 VPWR VGND sg13g2_decap_8
XFILLER_14_81 VPWR VGND sg13g2_decap_4
XFILLER_10_783 VPWR VGND sg13g2_decap_8
XFILLER_6_765 VPWR VGND sg13g2_decap_8
XFILLER_5_297 VPWR VGND sg13g2_fill_2
XFILLER_1_470 VPWR VGND sg13g2_decap_8
XFILLER_49_452 VPWR VGND sg13g2_decap_4
X_3000_ _1143_ net232 net613 VPWR VGND sg13g2_nand2_1
Xinput7 ui_in[5] net7 VPWR VGND sg13g2_buf_1
XFILLER_45_680 VPWR VGND sg13g2_decap_8
XFILLER_18_894 VPWR VGND sg13g2_fill_1
X_3902_ net945 net899 net599 _0414_ VPWR VGND sg13g2_mux2_1
XFILLER_33_853 VPWR VGND sg13g2_fill_1
X_3833_ _1740_ _1758_ _1759_ _1760_ VPWR VGND sg13g2_nor3_1
XFILLER_20_503 VPWR VGND sg13g2_fill_1
XFILLER_32_385 VPWR VGND sg13g2_fill_1
X_3764_ VGND VPWR _1709_ _1465_ _0589_ sg13g2_or2_1
X_2715_ _0971_ net521 net49 VPWR VGND sg13g2_nand2b_1
X_3695_ _1645_ VPWR _0345_ VGND _1663_ _1664_ sg13g2_o21ai_1
X_2646_ net913 net973 _0917_ VPWR VGND sg13g2_nor2_2
X_2577_ _0861_ VPWR _0015_ VGND _1919_ _0647_ sg13g2_o21ai_1
X_4316_ net692 VGND VPWR net461 u_usb_cdc.u_sie.delay_cnt_q\[2\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
X_4247_ net640 VGND VPWR net875 net36 clknet_leaf_3_clk sg13g2_dfrbpq_1
X_4178_ net647 VGND VPWR net181 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[14\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_27_113 VPWR VGND sg13g2_fill_1
X_3129_ _1221_ net223 net627 VPWR VGND sg13g2_nand2_1
XFILLER_24_820 VPWR VGND sg13g2_fill_2
XFILLER_23_352 VPWR VGND sg13g2_fill_1
XFILLER_3_724 VPWR VGND sg13g2_decap_8
XFILLER_47_912 VPWR VGND sg13g2_decap_8
Xfanout571 _1388_ net571 VPWR VGND sg13g2_buf_1
Xfanout582 _0869_ net582 VPWR VGND sg13g2_buf_8
Xfanout593 net596 net593 VPWR VGND sg13g2_buf_8
XFILLER_19_636 VPWR VGND sg13g2_fill_2
XFILLER_47_989 VPWR VGND sg13g2_decap_8
XFILLER_46_466 VPWR VGND sg13g2_fill_2
XFILLER_18_157 VPWR VGND sg13g2_fill_1
XFILLER_15_820 VPWR VGND sg13g2_decap_8
XFILLER_14_374 VPWR VGND sg13g2_decap_4
XFILLER_41_160 VPWR VGND sg13g2_fill_2
X_3480_ _1475_ net319 net289 VPWR VGND sg13g2_xnor2_1
X_2500_ VGND VPWR _0791_ _0796_ _0797_ _0739_ sg13g2_a21oi_1
XFILLER_6_573 VPWR VGND sg13g2_decap_8
X_2431_ _0728_ _0726_ _0729_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_1021 VPWR VGND sg13g2_decap_8
X_2362_ _0655_ _0661_ _0662_ VPWR VGND sg13g2_nor2_2
X_4101_ net651 VGND VPWR net94 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[21\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2293_ _0595_ _1904_ net597 VPWR VGND sg13g2_nand2_2
X_4032_ net689 VGND VPWR net851 u_usb_cdc.u_sie.out_toggle_q\[1\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
XFILLER_37_400 VPWR VGND sg13g2_decap_8
XFILLER_38_956 VPWR VGND sg13g2_decap_8
XFILLER_25_606 VPWR VGND sg13g2_fill_2
XFILLER_36_1003 VPWR VGND sg13g2_decap_8
X_3816_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[0\] u_usb_cdc.u_sie.u_phy_rx.cnt_q\[1\] net202
+ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[3\] _1747_ VPWR VGND sg13g2_and4_1
X_3747_ VGND VPWR _1696_ _0618_ _0577_ sg13g2_or2_1
X_3678_ VGND VPWR net802 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[14\]
+ _1648_ _1647_ sg13g2_a21oi_1
X_2629_ _0904_ net847 net595 VPWR VGND sg13g2_nand2_1
XFILLER_0_738 VPWR VGND sg13g2_decap_8
XFILLER_29_901 VPWR VGND sg13g2_decap_8
XFILLER_29_912 VPWR VGND sg13g2_fill_2
XFILLER_16_606 VPWR VGND sg13g2_fill_2
XFILLER_44_948 VPWR VGND sg13g2_decap_8
XFILLER_28_499 VPWR VGND sg13g2_decap_4
XFILLER_12_878 VPWR VGND sg13g2_decap_8
XFILLER_4_1023 VPWR VGND sg13g2_fill_2
XFILLER_4_1012 VPWR VGND sg13g2_decap_8
XFILLER_19_411 VPWR VGND sg13g2_decap_8
XFILLER_47_786 VPWR VGND sg13g2_decap_8
XFILLER_34_414 VPWR VGND sg13g2_decap_4
X_2980_ _1131_ VPWR _0163_ VGND _1912_ _1130_ sg13g2_o21ai_1
XFILLER_43_992 VPWR VGND sg13g2_decap_8
X_3601_ VGND VPWR net773 _1511_ _1575_ _0650_ sg13g2_a21oi_1
Xinput10 uio_in[0] net10 VPWR VGND sg13g2_buf_1
XFILLER_7_871 VPWR VGND sg13g2_decap_8
X_3532_ _1508_ _1507_ _0551_ VPWR VGND sg13g2_nand2b_1
X_3463_ net739 net1046 _1463_ VPWR VGND sg13g2_nor2b_1
X_2414_ _0656_ _0659_ net715 _0712_ VPWR VGND net617 sg13g2_nand4_1
X_3394_ net754 _1408_ _1417_ VPWR VGND sg13g2_nor2_1
X_2345_ net738 VPWR _0646_ VGND _0610_ _0622_ sg13g2_o21ai_1
X_2276_ _0578_ net946 net634 VPWR VGND sg13g2_nand2_2
X_4015_ net638 _1890_ net736 _1891_ VPWR VGND sg13g2_nand3_1
XFILLER_38_764 VPWR VGND sg13g2_fill_1
XFILLER_12_108 VPWR VGND sg13g2_fill_1
XFILLER_40_439 VPWR VGND sg13g2_fill_2
XFILLER_32_37 VPWR VGND sg13g2_decap_4
XFILLER_0_535 VPWR VGND sg13g2_decap_8
XFILLER_29_764 VPWR VGND sg13g2_decap_8
XFILLER_31_417 VPWR VGND sg13g2_decap_8
XFILLER_24_480 VPWR VGND sg13g2_fill_1
XFILLER_12_642 VPWR VGND sg13g2_decap_8
XFILLER_40_984 VPWR VGND sg13g2_decap_8
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_3_351 VPWR VGND sg13g2_fill_1
XFILLER_3_384 VPWR VGND sg13g2_decap_8
X_2130_ _0066_ _2007_ net623 _2000_ _1984_ VPWR VGND sg13g2_a22oi_1
XFILLER_47_550 VPWR VGND sg13g2_decap_8
X_2061_ VPWR _1940_ u_usb_cdc.u_sie.crc16_q\[13\] VGND sg13g2_inv_1
XFILLER_23_929 VPWR VGND sg13g2_fill_2
X_2963_ VGND VPWR _1122_ _1123_ _0621_ _0620_ sg13g2_a21oi_2
X_2894_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net452 _1098_ _0110_ VPWR VGND sg13g2_mux2_1
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
Xhold602 u_usb_cdc.u_ctrl_endp.rec_q\[0\] VPWR VGND net920 sg13g2_dlygate4sd3_1
Xhold635 u_usb_cdc.u_ctrl_endp.req_q\[3\] VPWR VGND net953 sg13g2_dlygate4sd3_1
Xhold624 u_usb_cdc.sie_out_data\[7\] VPWR VGND net942 sg13g2_dlygate4sd3_1
X_3515_ VGND VPWR net799 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[8\]
+ _1491_ _1490_ sg13g2_a21oi_1
Xhold613 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] VPWR VGND net931 sg13g2_dlygate4sd3_1
Xhold679 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[0\] VPWR VGND
+ net997 sg13g2_dlygate4sd3_1
Xhold646 u_usb_cdc.endp\[3\] VPWR VGND net964 sg13g2_dlygate4sd3_1
Xhold668 u_usb_cdc.u_sie.data_q\[0\] VPWR VGND net986 sg13g2_dlygate4sd3_1
Xhold657 u_usb_cdc.u_sie.phy_state_q\[11\] VPWR VGND net975 sg13g2_dlygate4sd3_1
X_3446_ _1451_ VPWR _0309_ VGND net719 net580 sg13g2_o21ai_1
X_3377_ _0673_ net617 _0752_ _1404_ VPWR VGND sg13g2_nor3_1
X_2328_ _0628_ VPWR _0629_ VGND u_usb_cdc.u_ctrl_endp.state_q\[1\] u_usb_cdc.u_ctrl_endp.state_q\[5\]
+ sg13g2_o21ai_1
X_2259_ net841 _0555_ _0557_ _0559_ _0561_ VPWR VGND sg13g2_nor4_1
XFILLER_38_572 VPWR VGND sg13g2_fill_2
XFILLER_43_47 VPWR VGND sg13g2_fill_2
XFILLER_22_962 VPWR VGND sg13g2_decap_4
XFILLER_5_638 VPWR VGND sg13g2_decap_8
XFILLER_0_332 VPWR VGND sg13g2_decap_8
XFILLER_1_855 VPWR VGND sg13g2_decap_8
XFILLER_49_837 VPWR VGND sg13g2_decap_8
XFILLER_44_586 VPWR VGND sg13g2_fill_1
XFILLER_31_225 VPWR VGND sg13g2_decap_8
XFILLER_40_781 VPWR VGND sg13g2_fill_1
XFILLER_9_966 VPWR VGND sg13g2_decap_8
X_3300_ _1356_ net805 _1357_ VPWR VGND sg13g2_xor2_1
X_4280_ net677 VGND VPWR _0282_ _0055_ clknet_leaf_47_clk sg13g2_dfrbpq_1
X_3231_ _1278_ _1299_ _1300_ _1301_ VPWR VGND sg13g2_nor3_1
X_3162_ _1238_ VPWR _0238_ VGND _1182_ _1229_ sg13g2_o21ai_1
XFILLER_27_509 VPWR VGND sg13g2_decap_4
X_2113_ net839 VPWR _1991_ VGND net706 _1988_ sg13g2_o21ai_1
X_3093_ _1201_ VPWR _0206_ VGND net717 net607 sg13g2_o21ai_1
XFILLER_35_520 VPWR VGND sg13g2_fill_1
X_2044_ VPWR _1923_ u_usb_cdc.u_sie.pid_q\[1\] VGND sg13g2_inv_1
XFILLER_35_597 VPWR VGND sg13g2_decap_8
X_3995_ _1877_ net327 net713 VPWR VGND sg13g2_nand2_1
XFILLER_31_770 VPWR VGND sg13g2_decap_8
X_2946_ net511 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net603 _0141_ VPWR VGND sg13g2_mux2_1
X_2877_ _1088_ VPWR _0102_ VGND net826 _1089_ sg13g2_o21ai_1
Xhold410 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[27\] VPWR VGND
+ net452 sg13g2_dlygate4sd3_1
Xhold421 _0145_ VPWR VGND net463 sg13g2_dlygate4sd3_1
Xhold454 _0245_ VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold443 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[2\] VPWR VGND net485 sg13g2_dlygate4sd3_1
Xhold432 _0114_ VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold476 u_usb_cdc.u_ctrl_endp.endp_q\[0\] VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold465 u_usb_cdc.u_sie.delay_cnt_q\[1\] VPWR VGND net507 sg13g2_dlygate4sd3_1
Xhold487 u_usb_cdc.u_sie.u_phy_rx.rx_valid_q VPWR VGND net529 sg13g2_dlygate4sd3_1
Xhold498 u_usb_cdc.u_sie.crc16_q\[9\] VPWR VGND net540 sg13g2_dlygate4sd3_1
X_3429_ _1443_ net951 _1424_ VPWR VGND sg13g2_nand2_1
XFILLER_38_391 VPWR VGND sg13g2_decap_8
XFILLER_41_501 VPWR VGND sg13g2_decap_8
XFILLER_26_597 VPWR VGND sg13g2_fill_1
XFILLER_13_247 VPWR VGND sg13g2_decap_8
XFILLER_16_1023 VPWR VGND sg13g2_decap_4
XFILLER_10_932 VPWR VGND sg13g2_decap_8
XFILLER_5_402 VPWR VGND sg13g2_decap_4
XFILLER_6_947 VPWR VGND sg13g2_decap_8
XFILLER_5_435 VPWR VGND sg13g2_decap_4
XFILLER_5_479 VPWR VGND sg13g2_decap_8
XFILLER_1_652 VPWR VGND sg13g2_decap_8
XFILLER_49_612 VPWR VGND sg13g2_fill_2
XFILLER_36_339 VPWR VGND sg13g2_fill_2
XFILLER_45_884 VPWR VGND sg13g2_decap_8
XFILLER_44_361 VPWR VGND sg13g2_fill_2
X_2800_ VGND VPWR u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ _1039_ _1041_ net997 sg13g2_a21oi_1
XFILLER_13_770 VPWR VGND sg13g2_decap_4
X_3780_ _1722_ _1720_ net485 net579 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[1\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_32_589 VPWR VGND sg13g2_decap_8
X_2731_ _0976_ VPWR _0979_ VGND _0977_ _0978_ sg13g2_o21ai_1
XFILLER_12_291 VPWR VGND sg13g2_decap_4
X_2662_ _0441_ VPWR _0931_ VGND _2008_ _2009_ sg13g2_o21ai_1
X_4401_ net728 VGND VPWR net359 u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_2593_ u_usb_cdc.u_sie.addr_q\[2\] u_usb_cdc.addr\[2\] _0874_ VPWR VGND sg13g2_xor2_1
X_4332_ net687 VGND VPWR net373 u_usb_cdc.u_sie.crc16_q\[11\] clknet_leaf_26_clk sg13g2_dfrbpq_1
X_4263_ net676 VGND VPWR _0265_ u_usb_cdc.u_ctrl_endp.endp_q\[2\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_1
X_3214_ _1286_ net806 _1279_ VPWR VGND sg13g2_nand2_1
X_4194_ net645 VGND VPWR net183 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[30\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_3145_ _1229_ net735 _1148_ VPWR VGND sg13g2_nand2_2
X_3076_ _1192_ VPWR _0198_ VGND net717 net609 sg13g2_o21ai_1
X_2027_ _1906_ net767 VPWR VGND sg13g2_inv_2
XFILLER_39_1001 VPWR VGND sg13g2_decap_8
X_3978_ _1865_ _1945_ u_usb_cdc.u_sie.phy_state_q\[4\] _1925_ net830 VPWR VGND sg13g2_a22oi_1
X_2929_ _1112_ net114 _1110_ VPWR VGND sg13g2_nand2_1
XFILLER_3_906 VPWR VGND sg13g2_decap_8
XFILLER_46_1005 VPWR VGND sg13g2_decap_8
Xhold240 u_usb_cdc.u_sie.u_phy_tx.data_q\[1\] VPWR VGND net282 sg13g2_dlygate4sd3_1
Xhold262 _0391_ VPWR VGND net304 sg13g2_dlygate4sd3_1
XFILLER_2_427 VPWR VGND sg13g2_decap_8
Xhold251 _0371_ VPWR VGND net293 sg13g2_dlygate4sd3_1
XFILLER_49_46 VPWR VGND sg13g2_decap_8
Xhold284 _0218_ VPWR VGND net326 sg13g2_dlygate4sd3_1
Xhold273 _0190_ VPWR VGND net315 sg13g2_dlygate4sd3_1
Xhold295 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[63\] VPWR VGND
+ net337 sg13g2_dlygate4sd3_1
XFILLER_49_68 VPWR VGND sg13g2_fill_2
XFILLER_49_57 VPWR VGND sg13g2_fill_2
Xfanout720 _1895_ net720 VPWR VGND sg13g2_buf_8
Xfanout742 net743 net742 VPWR VGND sg13g2_buf_8
Xfanout731 net732 net731 VPWR VGND sg13g2_buf_8
Xfanout753 net1014 net753 VPWR VGND sg13g2_buf_8
Xfanout775 net1030 net775 VPWR VGND sg13g2_buf_8
Xfanout764 net765 net764 VPWR VGND sg13g2_buf_8
Xfanout797 net804 net797 VPWR VGND sg13g2_buf_8
XFILLER_18_317 VPWR VGND sg13g2_decap_4
Xfanout786 net787 net786 VPWR VGND sg13g2_buf_8
XFILLER_33_309 VPWR VGND sg13g2_fill_2
XFILLER_14_501 VPWR VGND sg13g2_decap_8
XFILLER_26_383 VPWR VGND sg13g2_fill_2
XFILLER_27_884 VPWR VGND sg13g2_decap_4
XFILLER_14_556 VPWR VGND sg13g2_fill_1
XFILLER_10_740 VPWR VGND sg13g2_fill_1
XFILLER_6_744 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[6] net8 VPWR VGND sg13g2_buf_1
XFILLER_36_136 VPWR VGND sg13g2_decap_8
XFILLER_17_383 VPWR VGND sg13g2_fill_2
X_3901_ net940 net485 net599 _0413_ VPWR VGND sg13g2_mux2_1
X_3832_ VGND VPWR net172 _1753_ _1759_ net873 sg13g2_a21oi_1
XFILLER_9_560 VPWR VGND sg13g2_fill_2
X_3763_ net748 net750 _1707_ _1708_ VPWR VGND sg13g2_nor3_1
XFILLER_9_593 VPWR VGND sg13g2_decap_8
X_2714_ net49 _0970_ _0046_ VPWR VGND sg13g2_nor2_1
X_3694_ net597 VPWR _1664_ VGND net982 net624 sg13g2_o21ai_1
X_2645_ _0440_ _0913_ _0916_ VPWR VGND _0915_ sg13g2_nand3b_1
X_4315_ net692 VGND VPWR net509 u_usb_cdc.u_sie.delay_cnt_q\[1\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_2576_ u_usb_cdc.u_ctrl_endp.max_length_q\[6\] _0847_ _0848_ _0853_ _0861_ VPWR VGND
+ sg13g2_or4_1
X_4246_ net640 VGND VPWR net877 net35 clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4177_ net662 VGND VPWR net226 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[13\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
X_3128_ net820 _1964_ net737 _1220_ VPWR VGND _1183_ sg13g2_nand4_1
XFILLER_27_147 VPWR VGND sg13g2_fill_1
X_3059_ net822 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\]
+ _1183_ VPWR VGND sg13g2_and2_1
XFILLER_35_48 VPWR VGND sg13g2_fill_2
XFILLER_42_128 VPWR VGND sg13g2_fill_2
XFILLER_3_703 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_fill_1
XFILLER_2_246 VPWR VGND sg13g2_fill_2
Xfanout572 net573 net572 VPWR VGND sg13g2_buf_8
Xfanout583 _0637_ net583 VPWR VGND sg13g2_buf_8
XFILLER_18_125 VPWR VGND sg13g2_decap_4
Xfanout594 net596 net594 VPWR VGND sg13g2_buf_8
XFILLER_47_968 VPWR VGND sg13g2_decap_8
XFILLER_41_183 VPWR VGND sg13g2_fill_1
X_2430_ _1927_ u_usb_cdc.u_ctrl_endp.in_dir_q _1926_ _0728_ VPWR VGND sg13g2_nand3_1
XFILLER_29_1000 VPWR VGND sg13g2_decap_8
X_2361_ _0661_ _1915_ net716 VPWR VGND sg13g2_nand2_2
X_2292_ net747 net596 _0594_ VPWR VGND sg13g2_nor2_1
X_4100_ net669 VGND VPWR net62 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[20\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_49_250 VPWR VGND sg13g2_decap_8
X_4031_ net677 VGND VPWR net553 u_usb_cdc.u_ctrl_endp.req_q\[11\] clknet_leaf_50_clk
+ sg13g2_dfrbpq_1
XFILLER_38_935 VPWR VGND sg13g2_decap_8
XFILLER_49_294 VPWR VGND sg13g2_fill_1
XFILLER_37_456 VPWR VGND sg13g2_fill_2
XFILLER_25_629 VPWR VGND sg13g2_decap_4
XFILLER_37_478 VPWR VGND sg13g2_fill_2
XFILLER_18_692 VPWR VGND sg13g2_fill_1
XFILLER_24_128 VPWR VGND sg13g2_fill_2
XFILLER_24_139 VPWR VGND sg13g2_fill_2
XFILLER_33_673 VPWR VGND sg13g2_fill_1
XFILLER_21_846 VPWR VGND sg13g2_decap_8
X_3815_ _1745_ VPWR _0383_ VGND net202 _1746_ sg13g2_o21ai_1
XFILLER_21_857 VPWR VGND sg13g2_fill_2
XFILLER_21_868 VPWR VGND sg13g2_fill_2
X_3746_ _0581_ _0599_ _0999_ _1695_ VGND VPWR _1694_ sg13g2_nor4_2
X_3677_ net802 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[6\] _1647_
+ VPWR VGND sg13g2_nor2b_1
X_2628_ _0903_ VPWR _0026_ VGND _0616_ _0896_ sg13g2_o21ai_1
XFILLER_0_717 VPWR VGND sg13g2_decap_8
X_2559_ net864 net856 net523 u_usb_cdc.u_ctrl_endp.max_length_q\[3\] _0848_ VPWR VGND
+ sg13g2_or4_1
X_4229_ net639 VGND VPWR net146 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[65\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
XFILLER_29_979 VPWR VGND sg13g2_decap_8
XFILLER_44_927 VPWR VGND sg13g2_decap_8
XFILLER_15_117 VPWR VGND sg13g2_fill_1
XFILLER_28_489 VPWR VGND sg13g2_decap_4
XFILLER_23_172 VPWR VGND sg13g2_fill_1
XFILLER_3_566 VPWR VGND sg13g2_fill_1
XFILLER_19_423 VPWR VGND sg13g2_decap_4
XFILLER_47_765 VPWR VGND sg13g2_decap_8
XFILLER_46_242 VPWR VGND sg13g2_decap_8
XFILLER_34_437 VPWR VGND sg13g2_decap_8
XFILLER_34_448 VPWR VGND sg13g2_fill_1
XFILLER_43_971 VPWR VGND sg13g2_decap_8
XFILLER_15_651 VPWR VGND sg13g2_decap_8
XFILLER_30_654 VPWR VGND sg13g2_fill_1
X_3600_ net771 _1572_ _1573_ _1574_ VPWR VGND sg13g2_nor3_1
Xinput11 uio_in[2] net11 VPWR VGND sg13g2_buf_1
XFILLER_7_850 VPWR VGND sg13g2_decap_8
X_3531_ _1507_ _1429_ net780 VPWR VGND sg13g2_nand2b_1
X_3462_ net347 VPWR _0314_ VGND _1456_ _1462_ sg13g2_o21ai_1
X_2413_ net760 _0710_ _0711_ VPWR VGND sg13g2_nor2_1
X_3393_ net538 net567 _1416_ VPWR VGND sg13g2_nor2_1
X_2344_ _0610_ _0644_ net750 _0645_ VPWR VGND sg13g2_nand3_1
X_2275_ VPWR VGND net85 _0571_ net633 net165 _0577_ net634 sg13g2_a221oi_1
XFILLER_38_710 VPWR VGND sg13g2_decap_8
X_4014_ _1890_ net542 _1054_ VPWR VGND sg13g2_nand2_1
XFILLER_41_919 VPWR VGND sg13g2_decap_8
XFILLER_20_131 VPWR VGND sg13g2_fill_1
X_3729_ _1690_ VPWR _0353_ VGND _1901_ net598 sg13g2_o21ai_1
XFILLER_0_514 VPWR VGND sg13g2_decap_8
XFILLER_28_242 VPWR VGND sg13g2_fill_2
XFILLER_28_264 VPWR VGND sg13g2_fill_1
XFILLER_40_963 VPWR VGND sg13g2_decap_8
XFILLER_7_102 VPWR VGND sg13g2_decap_8
XFILLER_7_179 VPWR VGND sg13g2_fill_2
XFILLER_4_886 VPWR VGND sg13g2_decap_8
XFILLER_3_341 VPWR VGND sg13g2_fill_1
X_2060_ VPWR _1939_ u_usb_cdc.u_sie.crc16_q\[14\] VGND sg13g2_inv_1
XFILLER_47_90 VPWR VGND sg13g2_fill_1
XFILLER_23_919 VPWR VGND sg13g2_decap_4
X_2962_ _1122_ net739 net632 VPWR VGND sg13g2_nand2_1
XFILLER_33_1007 VPWR VGND sg13g2_decap_8
X_2893_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net426 _1098_ _0109_ VPWR VGND sg13g2_mux2_1
XFILLER_31_996 VPWR VGND sg13g2_decap_8
Xhold603 u_usb_cdc.u_ctrl_endp.req_q\[7\] VPWR VGND net921 sg13g2_dlygate4sd3_1
Xhold636 _0004_ VPWR VGND net954 sg13g2_dlygate4sd3_1
Xhold625 _0303_ VPWR VGND net943 sg13g2_dlygate4sd3_1
Xhold614 _0066_ VPWR VGND net932 sg13g2_dlygate4sd3_1
X_3514_ net799 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[0\] _1490_
+ VPWR VGND sg13g2_nor2b_1
X_3445_ _1451_ net200 net580 VPWR VGND sg13g2_nand2_1
Xhold647 _0306_ VPWR VGND net965 sg13g2_dlygate4sd3_1
Xhold669 u_usb_cdc.u_sie.u_phy_rx.state_q\[3\] VPWR VGND net987 sg13g2_dlygate4sd3_1
Xhold658 u_usb_cdc.u_sie.rx_valid VPWR VGND net976 sg13g2_dlygate4sd3_1
X_3376_ VGND VPWR _1900_ _1399_ _0287_ _1403_ sg13g2_a21oi_1
X_2327_ _0628_ u_usb_cdc.sie_in_req net634 VPWR VGND sg13g2_nand2_1
XFILLER_27_16 VPWR VGND sg13g2_decap_4
X_2258_ net841 _0557_ _0559_ _0560_ VPWR VGND sg13g2_nor3_1
XFILLER_26_713 VPWR VGND sg13g2_decap_8
XFILLER_27_38 VPWR VGND sg13g2_decap_8
X_2189_ _0491_ _0489_ _0490_ _0486_ _0485_ VPWR VGND sg13g2_a22oi_1
XFILLER_25_212 VPWR VGND sg13g2_decap_4
XFILLER_26_757 VPWR VGND sg13g2_fill_2
XFILLER_22_985 VPWR VGND sg13g2_decap_4
XFILLER_1_834 VPWR VGND sg13g2_decap_8
XFILLER_49_816 VPWR VGND sg13g2_decap_8
XFILLER_0_388 VPWR VGND sg13g2_decap_8
XFILLER_1_1016 VPWR VGND sg13g2_decap_8
XFILLER_1_1027 VPWR VGND sg13g2_fill_2
XFILLER_16_267 VPWR VGND sg13g2_decap_8
XFILLER_31_204 VPWR VGND sg13g2_fill_1
XFILLER_8_400 VPWR VGND sg13g2_fill_1
XFILLER_9_945 VPWR VGND sg13g2_decap_8
XFILLER_13_985 VPWR VGND sg13g2_decap_8
XFILLER_4_683 VPWR VGND sg13g2_decap_8
X_3230_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[26\] net815
+ _1300_ VPWR VGND sg13g2_nor2b_1
X_3161_ _1238_ net143 _1230_ VPWR VGND sg13g2_nand2_1
X_2112_ _1989_ net839 _1990_ VPWR VGND sg13g2_nor2b_1
XFILLER_48_882 VPWR VGND sg13g2_decap_8
X_3092_ _1201_ net141 net607 VPWR VGND sg13g2_nand2_1
X_2043_ VPWR _1922_ u_usb_cdc.u_sie.pid_q\[0\] VGND sg13g2_inv_1
X_3994_ net623 _1838_ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] _1876_ VPWR VGND _1875_
+ sg13g2_nand4_1
X_2945_ net434 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net603 _0140_ VPWR VGND sg13g2_mux2_1
X_2876_ _1089_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ _1082_ VPWR VGND sg13g2_nand2_1
Xhold411 _0110_ VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold400 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[1\] VPWR VGND
+ net442 sg13g2_dlygate4sd3_1
Xhold433 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[38\] VPWR VGND
+ net475 sg13g2_dlygate4sd3_1
Xhold422 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[66\] VPWR VGND
+ net464 sg13g2_dlygate4sd3_1
Xhold444 _1722_ VPWR VGND net486 sg13g2_dlygate4sd3_1
Xhold455 u_usb_cdc.u_sie.u_phy_rx.state_q\[2\] VPWR VGND net497 sg13g2_dlygate4sd3_1
Xhold466 _1470_ VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold477 u_usb_cdc.u_sie.u_phy_rx.rx_eop_q VPWR VGND net519 sg13g2_dlygate4sd3_1
Xhold499 _0501_ VPWR VGND net541 sg13g2_dlygate4sd3_1
Xhold488 _0045_ VPWR VGND net530 sg13g2_dlygate4sd3_1
X_3428_ _1439_ VPWR _0300_ VGND _1426_ _1442_ sg13g2_o21ai_1
X_3359_ net458 net571 _1394_ VPWR VGND sg13g2_nor2_1
XFILLER_39_860 VPWR VGND sg13g2_fill_1
XFILLER_13_237 VPWR VGND sg13g2_decap_4
XFILLER_16_1002 VPWR VGND sg13g2_decap_8
XFILLER_10_911 VPWR VGND sg13g2_decap_8
XFILLER_6_926 VPWR VGND sg13g2_decap_8
XFILLER_10_988 VPWR VGND sg13g2_decap_8
XFILLER_1_631 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_48_178 VPWR VGND sg13g2_decap_8
XFILLER_36_329 VPWR VGND sg13g2_fill_1
XFILLER_45_863 VPWR VGND sg13g2_decap_8
XFILLER_44_373 VPWR VGND sg13g2_fill_2
XFILLER_32_557 VPWR VGND sg13g2_fill_1
XFILLER_32_579 VPWR VGND sg13g2_fill_1
X_2730_ _0978_ u_usb_cdc.u_sie.phy_state_q\[9\] _0496_ VPWR VGND sg13g2_nand2_1
X_2661_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] VPWR _0930_ VGND _0444_ _0918_ sg13g2_o21ai_1
XFILLER_8_285 VPWR VGND sg13g2_fill_1
X_4400_ net724 VGND VPWR net879 u_usb_cdc.bus_reset clknet_leaf_37_clk sg13g2_dfrbpq_2
X_2592_ net837 net592 net746 _0873_ VPWR VGND sg13g2_nand3_1
X_4331_ net688 VGND VPWR _0333_ u_usb_cdc.u_sie.crc16_q\[10\] clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_5_981 VPWR VGND sg13g2_decap_8
XFILLER_5_52 VPWR VGND sg13g2_fill_2
X_4262_ net676 VGND VPWR _0264_ u_usb_cdc.u_ctrl_endp.endp_q\[1\] clknet_leaf_50_clk
+ sg13g2_dfrbpq_1
X_3213_ net805 _1284_ _1285_ VPWR VGND sg13g2_nor2_1
XFILLER_39_101 VPWR VGND sg13g2_fill_2
X_4193_ net663 VGND VPWR net205 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[29\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_1
X_3144_ _1228_ VPWR _0230_ VGND net717 net628 sg13g2_o21ai_1
X_3075_ _1192_ net201 net609 VPWR VGND sg13g2_nand2_1
XFILLER_36_830 VPWR VGND sg13g2_fill_2
X_2026_ VPWR _1905_ net884 VGND sg13g2_inv_1
XFILLER_23_535 VPWR VGND sg13g2_fill_1
XFILLER_24_28 VPWR VGND sg13g2_decap_8
X_3977_ _1864_ _1946_ net259 u_usb_cdc.u_sie.data_q\[7\] net834 VPWR VGND sg13g2_a22oi_1
XFILLER_11_708 VPWR VGND sg13g2_decap_4
X_2928_ _1111_ VPWR _0131_ VGND net707 _1083_ sg13g2_o21ai_1
X_2859_ _1075_ VPWR _0097_ VGND _1064_ _1076_ sg13g2_o21ai_1
XFILLER_2_406 VPWR VGND sg13g2_decap_8
Xhold241 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[21\] VPWR
+ VGND net283 sg13g2_dlygate4sd3_1
Xhold230 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[55\] VPWR
+ VGND net272 sg13g2_dlygate4sd3_1
Xhold252 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\] VPWR VGND net294 sg13g2_dlygate4sd3_1
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
Xhold263 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[15\] VPWR VGND net305 sg13g2_dlygate4sd3_1
Xhold296 _0146_ VPWR VGND net338 sg13g2_dlygate4sd3_1
Xhold285 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] VPWR VGND net327 sg13g2_dlygate4sd3_1
Xhold274 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[1\] VPWR VGND net316 sg13g2_dlygate4sd3_1
Xfanout721 _1894_ net721 VPWR VGND sg13g2_buf_8
Xfanout710 net712 net710 VPWR VGND sg13g2_buf_8
Xfanout732 net733 net732 VPWR VGND sg13g2_buf_8
Xfanout754 net996 net754 VPWR VGND sg13g2_buf_8
Xfanout743 net744 net743 VPWR VGND sg13g2_buf_8
Xfanout776 net777 net776 VPWR VGND sg13g2_buf_8
Xfanout765 net1052 net765 VPWR VGND sg13g2_buf_8
Xfanout798 net804 net798 VPWR VGND sg13g2_buf_8
Xfanout787 net1063 net787 VPWR VGND sg13g2_buf_8
XFILLER_42_800 VPWR VGND sg13g2_fill_1
XFILLER_10_796 VPWR VGND sg13g2_fill_2
XFILLER_6_723 VPWR VGND sg13g2_decap_8
XFILLER_5_222 VPWR VGND sg13g2_fill_2
XFILLER_5_266 VPWR VGND sg13g2_decap_4
XFILLER_2_984 VPWR VGND sg13g2_decap_8
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
XFILLER_49_498 VPWR VGND sg13g2_decap_8
Xinput9 ui_in[7] net9 VPWR VGND sg13g2_buf_1
XFILLER_37_638 VPWR VGND sg13g2_decap_4
XFILLER_17_395 VPWR VGND sg13g2_fill_2
X_3900_ net967 net531 net599 _0412_ VPWR VGND sg13g2_mux2_1
XFILLER_33_844 VPWR VGND sg13g2_decap_8
X_3831_ _1758_ net172 net873 _1753_ VPWR VGND sg13g2_and3_1
X_3762_ _1706_ _0908_ _1707_ VPWR VGND sg13g2_nor2b_1
X_2713_ _0970_ _0968_ _0969_ VPWR VGND sg13g2_nand2_1
X_3693_ VPWR VGND _1528_ _1489_ _1662_ net631 _1663_ _1659_ sg13g2_a221oi_1
X_2644_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] _0914_ _0915_ VPWR VGND sg13g2_and2_1
X_2575_ net947 VPWR _0014_ VGND _0680_ _0860_ sg13g2_o21ai_1
X_4314_ net691 VGND VPWR net1006 u_usb_cdc.u_sie.delay_cnt_q\[0\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_2
X_4245_ net640 VGND VPWR net898 net34 clknet_leaf_3_clk sg13g2_dfrbpq_1
X_4176_ net659 VGND VPWR net154 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[12\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3127_ VGND VPWR _1182_ net605 _0222_ _1219_ sg13g2_a21oi_1
XFILLER_28_638 VPWR VGND sg13g2_fill_1
X_3058_ VGND VPWR net612 _1182_ _0190_ _1181_ sg13g2_a21oi_1
XFILLER_24_822 VPWR VGND sg13g2_fill_1
XFILLER_24_877 VPWR VGND sg13g2_fill_1
XFILLER_11_516 VPWR VGND sg13g2_decap_4
XFILLER_23_387 VPWR VGND sg13g2_decap_4
XFILLER_13_1027 VPWR VGND sg13g2_fill_2
XFILLER_2_214 VPWR VGND sg13g2_decap_4
XFILLER_3_759 VPWR VGND sg13g2_decap_8
Xfanout573 _1484_ net573 VPWR VGND sg13g2_buf_8
Xfanout584 net585 net584 VPWR VGND sg13g2_buf_8
XFILLER_47_947 VPWR VGND sg13g2_decap_8
XFILLER_46_424 VPWR VGND sg13g2_fill_2
XFILLER_46_413 VPWR VGND sg13g2_fill_1
Xfanout595 net596 net595 VPWR VGND sg13g2_buf_8
XFILLER_42_630 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_53_clk clknet_3_1__leaf_clk clknet_leaf_53_clk VPWR VGND sg13g2_buf_8
X_2360_ net786 net785 _0660_ VPWR VGND sg13g2_nor2_1
XFILLER_2_781 VPWR VGND sg13g2_decap_8
X_2291_ _0593_ net743 _0590_ VPWR VGND sg13g2_nand2_1
XFILLER_49_240 VPWR VGND sg13g2_fill_1
X_4030_ net665 VGND VPWR net207 u_usb_cdc.u_ctrl_endp.req_q\[10\] clknet_leaf_49_clk
+ sg13g2_dfrbpq_1
XFILLER_25_608 VPWR VGND sg13g2_fill_1
XFILLER_46_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_44_clk clknet_3_4__leaf_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
XFILLER_24_118 VPWR VGND sg13g2_fill_2
X_3814_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[1\] net600 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[0\]
+ _1746_ VPWR VGND sg13g2_nand3_1
XFILLER_32_195 VPWR VGND sg13g2_fill_2
X_3745_ net836 _1693_ _1694_ VPWR VGND sg13g2_nor2_1
X_3676_ _1646_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[70\] net626
+ VPWR VGND sg13g2_nand2_1
X_2627_ _0903_ _0613_ _1904_ net593 net835 VPWR VGND sg13g2_a22oi_1
X_2558_ VGND VPWR _0847_ net854 net538 sg13g2_or2_1
X_2489_ _0781_ _0783_ _0785_ _0786_ VPWR VGND sg13g2_nor3_1
X_4228_ net639 VGND VPWR net119 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[64\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_28_424 VPWR VGND sg13g2_fill_2
XFILLER_44_906 VPWR VGND sg13g2_decap_8
X_4159_ net672 VGND VPWR _0162_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_29_958 VPWR VGND sg13g2_decap_8
XFILLER_43_438 VPWR VGND sg13g2_decap_8
XFILLER_24_641 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_35_clk clknet_3_6__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_11_313 VPWR VGND sg13g2_decap_8
XFILLER_3_545 VPWR VGND sg13g2_decap_8
XFILLER_3_534 VPWR VGND sg13g2_fill_2
XFILLER_47_744 VPWR VGND sg13g2_decap_8
XFILLER_19_457 VPWR VGND sg13g2_fill_2
XFILLER_28_991 VPWR VGND sg13g2_decap_8
XFILLER_43_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_3_6__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
Xinput12 usb_dn_rx_i net12 VPWR VGND sg13g2_buf_1
X_3530_ _0664_ _1505_ _1506_ VPWR VGND sg13g2_nor2_1
XFILLER_6_361 VPWR VGND sg13g2_fill_2
X_3461_ _1459_ VPWR _1462_ VGND _1932_ net345 sg13g2_o21ai_1
X_2412_ _0702_ _0707_ net720 _0710_ VPWR VGND sg13g2_nand3_1
X_3392_ VGND VPWR net568 _1415_ _0291_ _1414_ sg13g2_a21oi_1
X_2343_ VGND VPWR _0632_ _0643_ _0644_ net714 sg13g2_a21oi_1
X_4013_ net903 _1889_ _1123_ _0438_ VPWR VGND sg13g2_mux2_1
X_2274_ _0576_ net767 net706 VPWR VGND sg13g2_nand2_2
XFILLER_38_777 VPWR VGND sg13g2_decap_8
XFILLER_25_449 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_17_clk clknet_3_3__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_40_408 VPWR VGND sg13g2_fill_1
XFILLER_34_994 VPWR VGND sg13g2_decap_8
XFILLER_21_633 VPWR VGND sg13g2_decap_4
X_3728_ net590 _1683_ net985 _1690_ VPWR VGND sg13g2_nand3_1
X_3659_ _1629_ VPWR _1630_ VGND net800 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[37\]
+ sg13g2_o21ai_1
XFILLER_29_700 VPWR VGND sg13g2_fill_1
XFILLER_28_210 VPWR VGND sg13g2_fill_2
XFILLER_29_777 VPWR VGND sg13g2_fill_2
XFILLER_29_799 VPWR VGND sg13g2_fill_2
XFILLER_43_246 VPWR VGND sg13g2_fill_1
XFILLER_12_622 VPWR VGND sg13g2_decap_4
XFILLER_40_942 VPWR VGND sg13g2_decap_8
XFILLER_11_143 VPWR VGND sg13g2_decap_8
XFILLER_7_125 VPWR VGND sg13g2_decap_4
XFILLER_4_865 VPWR VGND sg13g2_decap_8
XFILLER_3_397 VPWR VGND sg13g2_fill_1
XFILLER_26_1015 VPWR VGND sg13g2_decap_8
XFILLER_47_596 VPWR VGND sg13g2_fill_2
XFILLER_47_585 VPWR VGND sg13g2_decap_4
XFILLER_35_758 VPWR VGND sg13g2_decap_4
X_2961_ net491 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ _1121_ _0154_ VPWR VGND sg13g2_mux2_1
XFILLER_8_30 VPWR VGND sg13g2_fill_1
XFILLER_31_975 VPWR VGND sg13g2_decap_8
X_2892_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net489 _1098_ _0108_ VPWR VGND sg13g2_mux2_1
Xhold604 _0008_ VPWR VGND net922 sg13g2_dlygate4sd3_1
Xhold626 u_usb_cdc.u_sie.rx_err VPWR VGND net944 sg13g2_dlygate4sd3_1
Xhold615 net28 VPWR VGND net933 sg13g2_dlygate4sd3_1
X_3513_ VGND VPWR _1489_ _1481_ net747 sg13g2_or2_1
X_3444_ _1450_ VPWR _0308_ VGND net718 net581 sg13g2_o21ai_1
Xclkbuf_leaf_6_clk clknet_3_1__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
Xhold659 _1800_ VPWR VGND net977 sg13g2_dlygate4sd3_1
Xhold637 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[0\] VPWR VGND
+ net955 sg13g2_dlygate4sd3_1
Xhold648 u_usb_cdc.u_sie.rx_data\[3\] VPWR VGND net966 sg13g2_dlygate4sd3_1
X_3375_ net993 _1399_ _1403_ VPWR VGND sg13g2_nor2_1
X_2326_ _0625_ VPWR _0627_ VGND _0610_ _0622_ sg13g2_o21ai_1
X_2257_ VGND VPWR _0559_ u_usb_cdc.u_ctrl_endp.state_q\[2\] u_usb_cdc.u_ctrl_endp.state_q\[1\]
+ sg13g2_or2_1
X_2188_ _0483_ u_usb_cdc.u_sie.data_q\[3\] _0490_ VPWR VGND sg13g2_xor2_1
XFILLER_25_224 VPWR VGND sg13g2_fill_2
XFILLER_26_747 VPWR VGND sg13g2_fill_1
XFILLER_21_496 VPWR VGND sg13g2_fill_2
XFILLER_4_106 VPWR VGND sg13g2_fill_2
XFILLER_49_1026 VPWR VGND sg13g2_fill_2
XFILLER_1_813 VPWR VGND sg13g2_decap_8
XFILLER_0_367 VPWR VGND sg13g2_decap_8
XFILLER_48_338 VPWR VGND sg13g2_fill_1
XFILLER_44_500 VPWR VGND sg13g2_fill_2
XFILLER_9_924 VPWR VGND sg13g2_decap_8
XFILLER_13_964 VPWR VGND sg13g2_decap_8
XFILLER_12_485 VPWR VGND sg13g2_fill_2
XFILLER_4_662 VPWR VGND sg13g2_decap_8
X_3160_ _1237_ VPWR _0237_ VGND _1180_ _1229_ sg13g2_o21ai_1
X_3091_ _1200_ VPWR _0205_ VGND _1901_ net607 sg13g2_o21ai_1
Xhold1 u_usb_cdc.u_sie.u_phy_rx.dn_q\[2\] VPWR VGND net43 sg13g2_dlygate4sd3_1
X_2111_ net706 _1988_ _1989_ VPWR VGND sg13g2_nor2_2
XFILLER_48_861 VPWR VGND sg13g2_decap_8
X_2042_ VPWR _1921_ net460 VGND sg13g2_inv_1
X_3993_ _1875_ _0586_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] VPWR VGND sg13g2_nand2b_1
X_2944_ net395 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net603 _0139_ VPWR VGND sg13g2_mux2_1
X_2875_ _1088_ net184 _1080_ VPWR VGND sg13g2_nand2_1
XFILLER_30_293 VPWR VGND sg13g2_decap_8
Xhold401 _0084_ VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold434 _0121_ VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold412 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[35\] VPWR VGND
+ net454 sg13g2_dlygate4sd3_1
Xhold423 _0149_ VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold445 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[60\] VPWR VGND
+ net487 sg13g2_dlygate4sd3_1
Xhold456 _0951_ VPWR VGND net498 sg13g2_dlygate4sd3_1
Xhold467 _0317_ VPWR VGND net509 sg13g2_dlygate4sd3_1
Xhold478 _0975_ VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold489 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[1\] VPWR VGND net531 sg13g2_dlygate4sd3_1
X_3427_ _1437_ net772 _1442_ VPWR VGND sg13g2_xor2_1
X_3358_ VGND VPWR _1899_ net571 _0279_ _1393_ sg13g2_a21oi_1
X_2309_ net634 _0609_ _0610_ VPWR VGND sg13g2_and2_1
XFILLER_46_809 VPWR VGND sg13g2_decap_8
X_3289_ net955 _1256_ _1352_ _0251_ VPWR VGND sg13g2_mux2_1
XFILLER_26_544 VPWR VGND sg13g2_decap_8
XFILLER_14_717 VPWR VGND sg13g2_decap_4
XFILLER_22_794 VPWR VGND sg13g2_fill_2
XFILLER_6_905 VPWR VGND sg13g2_decap_8
XFILLER_10_967 VPWR VGND sg13g2_decap_8
XFILLER_1_610 VPWR VGND sg13g2_decap_8
XFILLER_0_153 VPWR VGND sg13g2_fill_2
XFILLER_1_687 VPWR VGND sg13g2_decap_8
XFILLER_49_669 VPWR VGND sg13g2_decap_8
XFILLER_48_146 VPWR VGND sg13g2_fill_1
XFILLER_45_842 VPWR VGND sg13g2_decap_8
XFILLER_44_385 VPWR VGND sg13g2_fill_1
XFILLER_9_765 VPWR VGND sg13g2_decap_4
X_2660_ _0928_ VPWR _0002_ VGND _0741_ _0929_ sg13g2_o21ai_1
XFILLER_5_960 VPWR VGND sg13g2_decap_8
X_2591_ _0872_ net746 net592 VPWR VGND sg13g2_nand2_1
X_4330_ net687 VGND VPWR _0332_ u_usb_cdc.u_sie.crc16_q\[9\] clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_5_86 VPWR VGND sg13g2_fill_2
X_4261_ net676 VGND VPWR _0263_ u_usb_cdc.u_ctrl_endp.endp_q\[0\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
XFILLER_4_492 VPWR VGND sg13g2_fill_2
X_3212_ VPWR VGND _1280_ _1283_ _1279_ net808 _1284_ _1277_ sg13g2_a221oi_1
X_4192_ net661 VGND VPWR net177 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[28\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_1
X_3143_ _1228_ net161 net628 VPWR VGND sg13g2_nand2_1
X_3074_ _1191_ VPWR _0197_ VGND _1901_ net610 sg13g2_o21ai_1
X_2025_ net747 _1904_ VPWR VGND sg13g2_inv_4
XFILLER_36_864 VPWR VGND sg13g2_fill_1
X_3976_ VGND VPWR _1863_ _1696_ _1018_ sg13g2_or2_1
X_2927_ _1111_ net155 _1110_ VPWR VGND sg13g2_nand2_1
X_2858_ _1076_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2789_ net219 VPWR _0072_ VGND _0600_ _1031_ sg13g2_o21ai_1
Xhold220 _0063_ VPWR VGND net262 sg13g2_dlygate4sd3_1
Xhold242 _0188_ VPWR VGND net284 sg13g2_dlygate4sd3_1
Xhold231 _0222_ VPWR VGND net273 sg13g2_dlygate4sd3_1
Xhold253 _1792_ VPWR VGND net295 sg13g2_dlygate4sd3_1
Xhold264 u_usb_cdc.u_sie.crc16_q\[5\] VPWR VGND net306 sg13g2_dlygate4sd3_1
X_4459_ u_usb_cdc.configured_o net25 VPWR VGND sg13g2_buf_8
Xfanout700 net701 net700 VPWR VGND sg13g2_buf_8
Xhold286 _0433_ VPWR VGND net328 sg13g2_dlygate4sd3_1
Xhold275 _0434_ VPWR VGND net317 sg13g2_dlygate4sd3_1
Xhold297 u_usb_cdc.u_sie.in_byte_q\[3\] VPWR VGND net339 sg13g2_dlygate4sd3_1
Xfanout722 net724 net722 VPWR VGND sg13g2_buf_8
Xfanout733 net734 net733 VPWR VGND sg13g2_buf_8
Xfanout711 net713 net711 VPWR VGND sg13g2_buf_1
Xfanout755 net1016 net755 VPWR VGND sg13g2_buf_8
Xfanout744 net1049 net744 VPWR VGND sg13g2_buf_8
Xfanout766 net986 net766 VPWR VGND sg13g2_buf_8
Xfanout777 net778 net777 VPWR VGND sg13g2_buf_8
Xfanout788 net1048 net788 VPWR VGND sg13g2_buf_8
Xfanout799 net800 net799 VPWR VGND sg13g2_buf_8
XFILLER_41_300 VPWR VGND sg13g2_fill_2
XFILLER_26_385 VPWR VGND sg13g2_fill_1
XFILLER_41_366 VPWR VGND sg13g2_fill_2
XFILLER_6_779 VPWR VGND sg13g2_decap_8
XFILLER_30_61 VPWR VGND sg13g2_decap_4
XFILLER_30_94 VPWR VGND sg13g2_fill_2
XFILLER_2_963 VPWR VGND sg13g2_decap_8
XFILLER_1_484 VPWR VGND sg13g2_decap_8
XFILLER_49_477 VPWR VGND sg13g2_decap_8
XFILLER_18_853 VPWR VGND sg13g2_fill_1
XFILLER_45_694 VPWR VGND sg13g2_decap_8
XFILLER_17_385 VPWR VGND sg13g2_fill_1
X_3830_ VGND VPWR net172 _1755_ _0387_ _1757_ sg13g2_a21oi_1
XFILLER_13_580 VPWR VGND sg13g2_decap_8
X_3761_ _0529_ _0987_ _1706_ VPWR VGND sg13g2_nor2_1
X_2712_ _0969_ u_usb_cdc.u_sie.u_phy_rx.dp_q\[0\] net47 VPWR VGND sg13g2_xnor2_1
X_3692_ VGND VPWR _1662_ _1661_ _1636_ sg13g2_or2_1
X_2643_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\] u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[2\]
+ _0914_ VPWR VGND u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] sg13g2_nand3b_1
X_2574_ VGND VPWR _0681_ _0852_ _0860_ net584 sg13g2_a21oi_1
X_4313_ net686 VGND VPWR _0315_ u_usb_cdc.sie_in_req clknet_leaf_23_clk sg13g2_dfrbpq_2
X_4244_ net640 VGND VPWR net545 net33 clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4175_ net644 VGND VPWR net103 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[11\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3126_ net272 net605 _1219_ VPWR VGND sg13g2_nor2_1
XFILLER_43_609 VPWR VGND sg13g2_decap_8
X_3057_ _1182_ net751 _1135_ VPWR VGND sg13g2_nand2_2
X_3959_ _1848_ VPWR _1849_ VGND net274 net705 sg13g2_o21ai_1
XFILLER_13_1006 VPWR VGND sg13g2_decap_8
XFILLER_3_738 VPWR VGND sg13g2_decap_8
Xfanout574 _0693_ net574 VPWR VGND sg13g2_buf_8
XFILLER_47_926 VPWR VGND sg13g2_decap_8
Xfanout585 _0636_ net585 VPWR VGND sg13g2_buf_2
Xfanout596 _0593_ net596 VPWR VGND sg13g2_buf_8
XFILLER_46_436 VPWR VGND sg13g2_decap_4
XFILLER_26_160 VPWR VGND sg13g2_decap_8
XFILLER_26_171 VPWR VGND sg13g2_fill_2
XFILLER_2_760 VPWR VGND sg13g2_decap_8
X_2290_ net739 _0590_ _0592_ VPWR VGND sg13g2_and2_1
XFILLER_1_281 VPWR VGND sg13g2_fill_2
XFILLER_2_98 VPWR VGND sg13g2_decap_8
XFILLER_46_970 VPWR VGND sg13g2_decap_8
XFILLER_36_1017 VPWR VGND sg13g2_decap_8
X_3813_ net202 VPWR _1745_ VGND net712 _1742_ sg13g2_o21ai_1
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_369 VPWR VGND sg13g2_decap_8
X_3744_ VPWR _1693_ _1692_ VGND sg13g2_inv_1
X_3675_ _1645_ net985 net593 VPWR VGND sg13g2_nand2_1
X_2626_ _0902_ VPWR _0025_ VGND net208 _0872_ sg13g2_o21ai_1
X_2557_ net550 VPWR _0846_ VGND _0646_ _0845_ sg13g2_o21ai_1
X_2488_ _0709_ _0784_ _0785_ VPWR VGND sg13g2_nor2_1
X_4227_ net662 VGND VPWR _0230_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[63\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_28_403 VPWR VGND sg13g2_decap_8
X_4158_ net672 VGND VPWR _0161_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_43_417 VPWR VGND sg13g2_fill_2
X_3109_ _1210_ net112 _1202_ VPWR VGND sg13g2_nand2_1
X_4089_ net656 VGND VPWR net76 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[9\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_12_848 VPWR VGND sg13g2_fill_2
XFILLER_23_185 VPWR VGND sg13g2_fill_2
XFILLER_11_74 VPWR VGND sg13g2_fill_1
XFILLER_3_579 VPWR VGND sg13g2_decap_8
XFILLER_47_723 VPWR VGND sg13g2_decap_8
XFILLER_46_211 VPWR VGND sg13g2_fill_2
XFILLER_28_970 VPWR VGND sg13g2_decap_8
XFILLER_36_93 VPWR VGND sg13g2_decap_8
XFILLER_30_612 VPWR VGND sg13g2_fill_1
Xinput13 usb_dp_rx_i net13 VPWR VGND sg13g2_buf_1
XFILLER_30_689 VPWR VGND sg13g2_fill_2
XFILLER_11_881 VPWR VGND sg13g2_fill_1
XFILLER_7_885 VPWR VGND sg13g2_decap_8
XFILLER_6_351 VPWR VGND sg13g2_fill_1
X_3460_ _1461_ net346 _1456_ VPWR VGND sg13g2_nand2_1
X_2411_ net757 _0708_ _0709_ VPWR VGND sg13g2_nor2_1
X_3391_ net755 _1408_ _1415_ VPWR VGND sg13g2_nor2_1
X_2342_ _0556_ _0559_ _0643_ VPWR VGND sg13g2_nor2_1
X_4012_ _1041_ net828 _1054_ _1889_ VPWR VGND sg13g2_mux2_1
X_2273_ net767 net706 _0575_ VPWR VGND sg13g2_and2_1
XFILLER_37_222 VPWR VGND sg13g2_fill_2
XFILLER_34_973 VPWR VGND sg13g2_decap_8
XFILLER_21_689 VPWR VGND sg13g2_decap_8
X_3727_ _1689_ VPWR _0352_ VGND _1898_ net598 sg13g2_o21ai_1
XFILLER_10_1009 VPWR VGND sg13g2_decap_8
X_3658_ VGND VPWR net800 _1972_ _1629_ net793 sg13g2_a21oi_1
X_3589_ _1562_ VPWR _1563_ VGND net798 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[34\]
+ sg13g2_o21ai_1
X_2609_ _0890_ net766 _0889_ VPWR VGND sg13g2_nand2_2
XFILLER_48_509 VPWR VGND sg13g2_decap_8
XFILLER_0_549 VPWR VGND sg13g2_decap_8
XFILLER_44_715 VPWR VGND sg13g2_fill_2
XFILLER_44_737 VPWR VGND sg13g2_decap_8
XFILLER_40_921 VPWR VGND sg13g2_decap_8
XFILLER_19_1023 VPWR VGND sg13g2_decap_4
XFILLER_40_998 VPWR VGND sg13g2_decap_8
XFILLER_4_844 VPWR VGND sg13g2_decap_8
XFILLER_3_321 VPWR VGND sg13g2_fill_2
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_47_564 VPWR VGND sg13g2_decap_4
XFILLER_34_225 VPWR VGND sg13g2_fill_1
XFILLER_15_472 VPWR VGND sg13g2_fill_2
XFILLER_22_409 VPWR VGND sg13g2_decap_8
X_2960_ net469 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ _1121_ _0153_ VPWR VGND sg13g2_mux2_1
XFILLER_30_431 VPWR VGND sg13g2_decap_8
XFILLER_31_954 VPWR VGND sg13g2_decap_8
X_2891_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net418 _1098_ _0107_ VPWR VGND sg13g2_mux2_1
XFILLER_8_42 VPWR VGND sg13g2_fill_2
Xhold605 u_usb_cdc.u_sie.in_toggle_q\[1\] VPWR VGND net923 sg13g2_dlygate4sd3_1
Xhold616 _0365_ VPWR VGND net934 sg13g2_dlygate4sd3_1
Xhold627 u_usb_cdc.u_sie.rx_data\[2\] VPWR VGND net945 sg13g2_dlygate4sd3_1
X_3512_ net747 _1481_ _1488_ VPWR VGND sg13g2_nor2_1
X_3443_ _1450_ net213 net580 VPWR VGND sg13g2_nand2_1
Xhold638 _0251_ VPWR VGND net956 sg13g2_dlygate4sd3_1
Xhold649 u_usb_cdc.u_sie.rx_data\[0\] VPWR VGND net967 sg13g2_dlygate4sd3_1
X_3374_ VGND VPWR _1898_ _1399_ _0286_ _1402_ sg13g2_a21oi_1
X_2325_ VPWR _0626_ _0625_ VGND sg13g2_inv_1
X_2256_ VPWR _0558_ _0557_ VGND sg13g2_inv_1
X_2187_ _0489_ _0473_ _0488_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_759 VPWR VGND sg13g2_fill_1
XFILLER_13_409 VPWR VGND sg13g2_decap_8
XFILLER_22_921 VPWR VGND sg13g2_fill_1
XFILLER_21_431 VPWR VGND sg13g2_fill_2
XFILLER_33_280 VPWR VGND sg13g2_fill_2
XFILLER_33_291 VPWR VGND sg13g2_decap_8
XFILLER_21_486 VPWR VGND sg13g2_fill_2
XFILLER_49_1005 VPWR VGND sg13g2_decap_8
XFILLER_0_346 VPWR VGND sg13g2_decap_8
XFILLER_1_869 VPWR VGND sg13g2_decap_8
XFILLER_17_73 VPWR VGND sg13g2_decap_4
XFILLER_9_903 VPWR VGND sg13g2_decap_8
XFILLER_13_943 VPWR VGND sg13g2_decap_8
XFILLER_32_1020 VPWR VGND sg13g2_decap_8
XFILLER_8_479 VPWR VGND sg13g2_decap_8
XFILLER_8_468 VPWR VGND sg13g2_fill_1
XFILLER_4_641 VPWR VGND sg13g2_decap_8
XFILLER_3_195 VPWR VGND sg13g2_decap_4
X_3090_ _1200_ net139 net607 VPWR VGND sg13g2_nand2_1
Xhold2 u_usb_cdc.u_sie.u_phy_rx.dp_q\[2\] VPWR VGND net44 sg13g2_dlygate4sd3_1
X_2110_ net767 u_usb_cdc.endp\[3\] u_usb_cdc.endp\[2\] _1988_ VPWR VGND sg13g2_nor3_1
XFILLER_48_840 VPWR VGND sg13g2_decap_8
X_2041_ VPWR _1920_ net1003 VGND sg13g2_inv_1
XFILLER_35_545 VPWR VGND sg13g2_decap_4
X_3992_ _1874_ VPWR _0432_ VGND net741 _1980_ sg13g2_o21ai_1
XFILLER_23_729 VPWR VGND sg13g2_fill_2
X_2943_ _1043_ net615 _1119_ VPWR VGND sg13g2_nor2_2
X_2874_ _1086_ VPWR _0101_ VGND net826 _1087_ sg13g2_o21ai_1
XFILLER_30_272 VPWR VGND sg13g2_fill_2
XFILLER_31_784 VPWR VGND sg13g2_decap_4
Xhold402 u_usb_cdc.u_sie.crc16_q\[10\] VPWR VGND net444 sg13g2_dlygate4sd3_1
XFILLER_8_980 VPWR VGND sg13g2_decap_8
Xhold413 _0118_ VPWR VGND net455 sg13g2_dlygate4sd3_1
Xhold424 u_usb_cdc.u_sie.u_phy_tx.data_q\[4\] VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold435 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[67\] VPWR VGND
+ net477 sg13g2_dlygate4sd3_1
Xhold468 u_usb_cdc.u_ctrl_endp.addr_dd\[3\] VPWR VGND net510 sg13g2_dlygate4sd3_1
Xhold457 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[53\] VPWR
+ VGND net499 sg13g2_dlygate4sd3_1
Xhold446 _0143_ VPWR VGND net488 sg13g2_dlygate4sd3_1
Xhold479 u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[1\] VPWR VGND net521 sg13g2_dlygate4sd3_1
X_3426_ _1434_ _1440_ _1441_ VPWR VGND sg13g2_nor2_1
X_3357_ net384 net570 _1393_ VPWR VGND sg13g2_nor2_1
X_2308_ _0609_ _0608_ _0605_ VPWR VGND sg13g2_nand2b_1
X_3288_ net749 _0605_ _1239_ _1352_ VPWR VGND sg13g2_nor3_2
X_2239_ _0541_ net785 VPWR VGND net780 sg13g2_nand2b_2
XFILLER_26_534 VPWR VGND sg13g2_decap_4
XFILLER_22_762 VPWR VGND sg13g2_decap_4
XFILLER_10_946 VPWR VGND sg13g2_decap_8
XFILLER_1_666 VPWR VGND sg13g2_decap_8
XFILLER_49_648 VPWR VGND sg13g2_decap_8
XFILLER_23_1008 VPWR VGND sg13g2_fill_2
XFILLER_23_1019 VPWR VGND sg13g2_decap_8
XFILLER_45_821 VPWR VGND sg13g2_decap_8
XFILLER_45_898 VPWR VGND sg13g2_decap_8
XFILLER_32_504 VPWR VGND sg13g2_decap_8
XFILLER_32_548 VPWR VGND sg13g2_decap_8
XFILLER_44_93 VPWR VGND sg13g2_fill_2
XFILLER_9_733 VPWR VGND sg13g2_decap_4
XFILLER_8_276 VPWR VGND sg13g2_decap_8
X_2590_ _0871_ net413 net595 VPWR VGND sg13g2_nand2_1
XFILLER_5_54 VPWR VGND sg13g2_fill_1
XFILLER_5_98 VPWR VGND sg13g2_fill_2
X_4260_ net673 VGND VPWR _0262_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_2
X_4191_ net644 VGND VPWR _0194_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[27\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3211_ _1278_ _1281_ _1282_ _1283_ VPWR VGND sg13g2_nor3_1
X_3142_ _1227_ VPWR _0229_ VGND _1901_ net629 sg13g2_o21ai_1
X_3073_ _1191_ net182 net610 VPWR VGND sg13g2_nand2_1
X_2024_ VPWR _1903_ net833 VGND sg13g2_inv_1
XFILLER_39_1015 VPWR VGND sg13g2_decap_8
X_3975_ VPWR _0427_ net401 VGND sg13g2_inv_1
X_2926_ _1057_ _1079_ net824 _1110_ VPWR VGND sg13g2_nand3_1
X_2857_ _1075_ net151 _1059_ VPWR VGND sg13g2_nand2_1
Xhold210 u_usb_cdc.u_sie.addr_q\[1\] VPWR VGND net252 sg13g2_dlygate4sd3_1
X_2788_ VGND VPWR net761 _0870_ _1031_ _1029_ sg13g2_a21oi_1
Xhold243 u_usb_cdc.u_sie.crc16_q\[4\] VPWR VGND net285 sg13g2_dlygate4sd3_1
Xhold232 u_usb_cdc.u_sie.u_phy_tx.data_q\[5\] VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold221 u_usb_cdc.u_sie.u_phy_rx.rx_err_q VPWR VGND net263 sg13g2_dlygate4sd3_1
XFILLER_46_1019 VPWR VGND sg13g2_decap_8
Xhold265 _0336_ VPWR VGND net307 sg13g2_dlygate4sd3_1
Xhold276 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[0\] VPWR VGND net318 sg13g2_dlygate4sd3_1
Xhold287 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[54\] VPWR
+ VGND net329 sg13g2_dlygate4sd3_1
X_4458_ u_usb_cdc.dp_pu_o net24 VPWR VGND sg13g2_buf_1
Xhold254 _0400_ VPWR VGND net296 sg13g2_dlygate4sd3_1
Xhold298 _0322_ VPWR VGND net340 sg13g2_dlygate4sd3_1
Xfanout723 net724 net723 VPWR VGND sg13g2_buf_8
Xfanout701 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.rstn net701 VPWR VGND sg13g2_buf_8
Xfanout712 net713 net712 VPWR VGND sg13g2_buf_8
X_3409_ _1428_ net785 _1424_ VPWR VGND sg13g2_nand2_1
X_4389_ net723 VGND VPWR net304 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[10\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
Xfanout756 net1062 net756 VPWR VGND sg13g2_buf_8
Xfanout745 net746 net745 VPWR VGND sg13g2_buf_8
Xfanout767 u_usb_cdc.endp\[0\] net767 VPWR VGND sg13g2_buf_8
Xfanout734 net1036 net734 VPWR VGND sg13g2_buf_8
Xfanout789 net790 net789 VPWR VGND sg13g2_buf_8
Xfanout778 net779 net778 VPWR VGND sg13g2_buf_8
XFILLER_38_180 VPWR VGND sg13g2_fill_2
XFILLER_27_876 VPWR VGND sg13g2_decap_4
XFILLER_14_515 VPWR VGND sg13g2_fill_2
XFILLER_14_537 VPWR VGND sg13g2_decap_4
XFILLER_26_375 VPWR VGND sg13g2_decap_4
XFILLER_27_898 VPWR VGND sg13g2_decap_4
XFILLER_41_389 VPWR VGND sg13g2_decap_4
XFILLER_14_85 VPWR VGND sg13g2_fill_2
XFILLER_22_592 VPWR VGND sg13g2_fill_1
XFILLER_6_758 VPWR VGND sg13g2_decap_8
XFILLER_5_224 VPWR VGND sg13g2_fill_1
XFILLER_2_942 VPWR VGND sg13g2_decap_8
XFILLER_49_423 VPWR VGND sg13g2_fill_1
XFILLER_49_412 VPWR VGND sg13g2_fill_2
XFILLER_1_463 VPWR VGND sg13g2_decap_8
XFILLER_49_456 VPWR VGND sg13g2_fill_1
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_18_810 VPWR VGND sg13g2_fill_2
X_3760_ net1018 _1705_ _1695_ _0369_ VPWR VGND sg13g2_mux2_1
X_2711_ _0968_ net386 net46 VPWR VGND sg13g2_xnor2_1
X_3691_ _0544_ _1516_ _1617_ _1660_ _1661_ VPWR VGND sg13g2_nor4_1
X_2642_ _0446_ _0911_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[7\] _0913_ VPWR VGND
+ _0912_ sg13g2_nand4_1
X_2573_ _0859_ net946 _0854_ VPWR VGND sg13g2_nand2b_1
X_4312_ net734 VGND VPWR net348 u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\] clknet_leaf_48_clk
+ sg13g2_dfrbpq_2
X_4243_ net640 VGND VPWR net560 net32 clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4174_ net645 VGND VPWR net123 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[10\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3125_ VGND VPWR _1180_ net605 _0221_ _1218_ sg13g2_a21oi_1
X_3056_ net314 net612 _1181_ VPWR VGND sg13g2_nor2_1
XFILLER_27_128 VPWR VGND sg13g2_fill_2
XFILLER_23_312 VPWR VGND sg13g2_decap_8
XFILLER_23_345 VPWR VGND sg13g2_decap_8
XFILLER_35_194 VPWR VGND sg13g2_decap_8
X_3958_ _1847_ _1808_ _1807_ _1848_ VPWR VGND sg13g2_a21o_1
X_2909_ _1057_ _1061_ net824 _1101_ VPWR VGND sg13g2_nand3_1
X_3889_ _1798_ VPWR _1799_ VGND u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] net346 sg13g2_o21ai_1
XFILLER_3_717 VPWR VGND sg13g2_decap_8
XFILLER_2_205 VPWR VGND sg13g2_decap_4
XFILLER_47_905 VPWR VGND sg13g2_decap_8
Xfanout575 net577 net575 VPWR VGND sg13g2_buf_8
Xfanout586 net587 net586 VPWR VGND sg13g2_buf_8
Xfanout597 _0592_ net597 VPWR VGND sg13g2_buf_8
XFILLER_46_426 VPWR VGND sg13g2_fill_1
XFILLER_14_312 VPWR VGND sg13g2_fill_2
XFILLER_14_323 VPWR VGND sg13g2_fill_2
XFILLER_14_367 VPWR VGND sg13g2_decap_8
XFILLER_14_378 VPWR VGND sg13g2_fill_2
XFILLER_23_890 VPWR VGND sg13g2_fill_2
XFILLER_10_540 VPWR VGND sg13g2_decap_8
XFILLER_6_544 VPWR VGND sg13g2_fill_2
XFILLER_29_1014 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_fill_1
XFILLER_49_264 VPWR VGND sg13g2_decap_4
XFILLER_38_949 VPWR VGND sg13g2_decap_8
X_3812_ _1743_ _1744_ _0382_ VPWR VGND sg13g2_nor2_1
XFILLER_33_687 VPWR VGND sg13g2_fill_1
X_3743_ net833 net840 _1692_ VPWR VGND sg13g2_nor2_2
X_3674_ _1626_ VPWR _0344_ VGND net593 _1644_ sg13g2_o21ai_1
X_2625_ _0902_ net837 net595 VPWR VGND sg13g2_nand2_1
X_2556_ _0844_ _0628_ _0845_ VPWR VGND sg13g2_nor2b_1
X_2487_ net842 _0688_ net738 _0784_ VPWR VGND sg13g2_nand3_1
X_4226_ net646 VGND VPWR net129 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[62\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4157_ net672 VGND VPWR _0160_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[1\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_2
X_3108_ _1209_ VPWR _0213_ VGND net708 _1163_ sg13g2_o21ai_1
XFILLER_28_448 VPWR VGND sg13g2_decap_4
X_4088_ net655 VGND VPWR net96 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[8\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
X_3039_ _1170_ net759 net630 VPWR VGND sg13g2_nand2_2
XFILLER_37_982 VPWR VGND sg13g2_decap_8
XFILLER_23_131 VPWR VGND sg13g2_decap_4
XFILLER_12_827 VPWR VGND sg13g2_fill_2
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1005 VPWR VGND sg13g2_decap_8
XFILLER_19_404 VPWR VGND sg13g2_decap_8
XFILLER_47_779 VPWR VGND sg13g2_decap_8
XFILLER_19_459 VPWR VGND sg13g2_fill_1
XFILLER_34_407 VPWR VGND sg13g2_decap_8
XFILLER_46_278 VPWR VGND sg13g2_fill_2
XFILLER_43_985 VPWR VGND sg13g2_decap_8
XFILLER_14_142 VPWR VGND sg13g2_fill_2
XFILLER_15_665 VPWR VGND sg13g2_decap_4
XFILLER_15_687 VPWR VGND sg13g2_decap_4
XFILLER_30_635 VPWR VGND sg13g2_decap_4
XFILLER_7_831 VPWR VGND sg13g2_decap_4
XFILLER_7_864 VPWR VGND sg13g2_decap_8
X_2410_ _0708_ _0702_ _0707_ VPWR VGND sg13g2_nand2_1
X_3390_ net916 net567 _1414_ VPWR VGND sg13g2_nor2_1
X_2341_ net535 _0641_ _0642_ VPWR VGND u_usb_cdc.u_ctrl_endp.state_q\[3\] sg13g2_nand3b_1
X_2272_ _1906_ _1985_ _0574_ VPWR VGND sg13g2_nor2_1
X_4011_ _1888_ VPWR _0437_ VGND _1910_ _1887_ sg13g2_o21ai_1
XFILLER_19_971 VPWR VGND sg13g2_fill_2
XFILLER_34_952 VPWR VGND sg13g2_decap_8
XFILLER_33_440 VPWR VGND sg13g2_fill_1
X_3726_ net591 _1683_ net995 _1689_ VPWR VGND sg13g2_nand3_1
X_3657_ net797 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[5\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[13\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[21\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[29\]
+ net791 _1628_ VPWR VGND sg13g2_mux4_1
X_3588_ VGND VPWR net800 _1969_ _1562_ net791 sg13g2_a21oi_1
X_2608_ _0885_ _0886_ _0887_ _0889_ VGND VPWR _0888_ sg13g2_nor4_2
XFILLER_0_528 VPWR VGND sg13g2_decap_8
X_2539_ _0691_ _0712_ _0678_ _0832_ VPWR VGND sg13g2_nand3_1
X_4209_ net662 VGND VPWR net109 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[45\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_29_779 VPWR VGND sg13g2_fill_1
XFILLER_44_749 VPWR VGND sg13g2_decap_4
XFILLER_40_900 VPWR VGND sg13g2_decap_8
XFILLER_40_977 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
XFILLER_3_377 VPWR VGND sg13g2_decap_8
XFILLER_47_543 VPWR VGND sg13g2_decap_8
X_2890_ VGND VPWR _1098_ net616 _1043_ sg13g2_or2_1
XFILLER_15_495 VPWR VGND sg13g2_fill_1
XFILLER_30_487 VPWR VGND sg13g2_fill_2
Xhold617 u_usb_cdc.u_sie.u_phy_rx.rx_en_q VPWR VGND net935 sg13g2_dlygate4sd3_1
Xhold606 _1021_ VPWR VGND net924 sg13g2_dlygate4sd3_1
X_3511_ _1487_ net766 net594 VPWR VGND sg13g2_nand2_1
X_3442_ _1449_ VPWR _0307_ VGND _1895_ net580 sg13g2_o21ai_1
Xhold628 u_usb_cdc.ctrl_stall VPWR VGND net946 sg13g2_dlygate4sd3_1
Xhold639 u_usb_cdc.u_sie.pid_q\[1\] VPWR VGND net957 sg13g2_dlygate4sd3_1
X_3373_ net884 _1399_ _1402_ VPWR VGND sg13g2_nor2_1
X_2324_ _0610_ VPWR _0625_ VGND net749 _0623_ sg13g2_o21ai_1
XFILLER_26_0 VPWR VGND sg13g2_fill_2
X_2255_ u_usb_cdc.u_ctrl_endp.state_q\[1\] u_usb_cdc.ctrl_stall u_usb_cdc.u_ctrl_endp.state_q\[5\]
+ _0556_ _0557_ VPWR VGND sg13g2_or4_1
X_2186_ _0488_ u_usb_cdc.sie_out_data\[3\] net766 VPWR VGND sg13g2_xnor2_1
XFILLER_38_543 VPWR VGND sg13g2_decap_4
XFILLER_38_565 VPWR VGND sg13g2_decap_8
XFILLER_21_410 VPWR VGND sg13g2_decap_8
XFILLER_21_421 VPWR VGND sg13g2_fill_1
XFILLER_22_944 VPWR VGND sg13g2_fill_2
XFILLER_22_955 VPWR VGND sg13g2_decap_8
XFILLER_4_108 VPWR VGND sg13g2_fill_1
X_3709_ VGND VPWR _1666_ _1677_ _1678_ _0576_ sg13g2_a21oi_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_848 VPWR VGND sg13g2_decap_8
XFILLER_16_226 VPWR VGND sg13g2_decap_4
XFILLER_12_410 VPWR VGND sg13g2_decap_8
XFILLER_13_922 VPWR VGND sg13g2_decap_8
XFILLER_31_218 VPWR VGND sg13g2_decap_8
XFILLER_40_741 VPWR VGND sg13g2_fill_2
XFILLER_24_292 VPWR VGND sg13g2_decap_8
XFILLER_9_959 VPWR VGND sg13g2_decap_8
XFILLER_13_999 VPWR VGND sg13g2_decap_8
XFILLER_3_163 VPWR VGND sg13g2_fill_1
XFILLER_4_697 VPWR VGND sg13g2_decap_8
XFILLER_0_892 VPWR VGND sg13g2_decap_8
Xhold3 u_usb_cdc.rstn_sq\[1\] VPWR VGND net45 sg13g2_dlygate4sd3_1
X_2040_ VPWR _1919_ net866 VGND sg13g2_inv_1
XFILLER_48_896 VPWR VGND sg13g2_decap_8
X_3991_ _0440_ _0917_ net741 _1874_ VPWR VGND sg13g2_nand3_1
X_2942_ _1118_ VPWR _0138_ VGND _1965_ _1097_ sg13g2_o21ai_1
X_2873_ _1087_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ _1082_ VPWR VGND sg13g2_nand2_1
Xhold414 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[30\] VPWR VGND
+ net456 sg13g2_dlygate4sd3_1
Xhold403 _0523_ VPWR VGND net445 sg13g2_dlygate4sd3_1
Xhold436 _0150_ VPWR VGND net478 sg13g2_dlygate4sd3_1
Xhold425 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[36\] VPWR VGND
+ net467 sg13g2_dlygate4sd3_1
Xhold469 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[58\] VPWR VGND
+ net511 sg13g2_dlygate4sd3_1
Xhold458 _1217_ VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold447 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[25\] VPWR VGND
+ net489 sg13g2_dlygate4sd3_1
X_3425_ _1440_ net775 net772 VPWR VGND sg13g2_nand2_1
X_3356_ VGND VPWR net719 net570 _0278_ _1392_ sg13g2_a21oi_1
X_3287_ _0250_ _1351_ _1350_ VPWR VGND sg13g2_nand2b_1
X_2307_ u_usb_cdc.u_sie.delay_cnt_q\[1\] u_usb_cdc.u_sie.delay_cnt_q\[0\] u_usb_cdc.u_sie.delay_cnt_q\[2\]
+ _0608_ VPWR VGND _0607_ sg13g2_nand4_1
X_2238_ _0534_ _0536_ _0537_ _0538_ _0540_ VPWR VGND sg13g2_nor4_1
XFILLER_39_852 VPWR VGND sg13g2_fill_2
XFILLER_39_896 VPWR VGND sg13g2_decap_8
X_2169_ _0471_ net756 net751 VPWR VGND sg13g2_xnor2_1
XFILLER_13_207 VPWR VGND sg13g2_fill_2
XFILLER_16_1016 VPWR VGND sg13g2_decap_8
XFILLER_10_925 VPWR VGND sg13g2_decap_8
XFILLER_16_1027 VPWR VGND sg13g2_fill_2
XFILLER_5_406 VPWR VGND sg13g2_fill_2
XFILLER_0_111 VPWR VGND sg13g2_fill_1
XFILLER_0_133 VPWR VGND sg13g2_fill_2
XFILLER_1_645 VPWR VGND sg13g2_decap_8
XFILLER_17_513 VPWR VGND sg13g2_decap_4
XFILLER_28_84 VPWR VGND sg13g2_decap_4
XFILLER_29_340 VPWR VGND sg13g2_fill_2
XFILLER_45_877 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_fill_1
XFILLER_13_763 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_fill_1
XFILLER_40_560 VPWR VGND sg13g2_fill_2
XFILLER_5_995 VPWR VGND sg13g2_decap_8
X_4190_ net661 VGND VPWR _0193_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[26\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3210_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[24\] net815
+ _1282_ VPWR VGND sg13g2_nor2b_1
X_3141_ _1227_ net128 net629 VPWR VGND sg13g2_nand2_1
X_3072_ _1190_ VPWR _0196_ VGND _1898_ net608 sg13g2_o21ai_1
X_2023_ VPWR _1902_ net745 VGND sg13g2_inv_1
X_3974_ _1862_ _1824_ _1861_ net621 net400 VPWR VGND sg13g2_a22oi_1
X_2925_ _1109_ VPWR _0130_ VGND _1078_ _1099_ sg13g2_o21ai_1
X_2856_ _1073_ VPWR _0096_ VGND net616 _1074_ sg13g2_o21ai_1
Xhold211 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[13\] VPWR VGND
+ net253 sg13g2_dlygate4sd3_1
Xhold200 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[32\] VPWR
+ VGND net242 sg13g2_dlygate4sd3_1
X_2787_ _1030_ net218 _0600_ VPWR VGND sg13g2_nand2_1
Xhold244 _0335_ VPWR VGND net286 sg13g2_dlygate4sd3_1
Xhold233 _0426_ VPWR VGND net275 sg13g2_dlygate4sd3_1
Xhold222 _0974_ VPWR VGND net264 sg13g2_dlygate4sd3_1
Xhold277 u_usb_cdc.u_sie.in_byte_q\[1\] VPWR VGND net319 sg13g2_dlygate4sd3_1
Xhold255 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[14\] VPWR VGND net297 sg13g2_dlygate4sd3_1
X_4457_ u_usb_cdc.in_ready_o[0] net23 VPWR VGND sg13g2_buf_1
Xhold266 _0054_ VPWR VGND net308 sg13g2_dlygate4sd3_1
XFILLER_49_39 VPWR VGND sg13g2_decap_8
Xhold299 u_usb_cdc.u_ctrl_endp.endp_q\[2\] VPWR VGND net341 sg13g2_dlygate4sd3_1
Xhold288 _0221_ VPWR VGND net330 sg13g2_dlygate4sd3_1
Xfanout724 net733 net724 VPWR VGND sg13g2_buf_8
Xfanout713 net714 net713 VPWR VGND sg13g2_buf_8
X_3408_ VGND VPWR _1915_ _1426_ _0295_ _1427_ sg13g2_a21oi_1
Xfanout702 _0954_ net702 VPWR VGND sg13g2_buf_8
Xfanout757 net758 net757 VPWR VGND sg13g2_buf_8
X_4388_ net723 VGND VPWR net394 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[9\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xfanout735 net737 net735 VPWR VGND sg13g2_buf_8
Xfanout746 net976 net746 VPWR VGND sg13g2_buf_8
X_3339_ _1385_ VPWR _0268_ VGND _1954_ _1384_ sg13g2_o21ai_1
Xfanout768 net769 net768 VPWR VGND sg13g2_buf_8
Xfanout779 net1061 net779 VPWR VGND sg13g2_buf_8
XFILLER_45_129 VPWR VGND sg13g2_decap_8
XFILLER_27_888 VPWR VGND sg13g2_fill_2
XFILLER_41_302 VPWR VGND sg13g2_fill_1
XFILLER_14_549 VPWR VGND sg13g2_decap_8
XFILLER_6_737 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_8
XFILLER_1_442 VPWR VGND sg13g2_decap_8
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
XFILLER_2_998 VPWR VGND sg13g2_decap_8
XFILLER_44_140 VPWR VGND sg13g2_fill_2
XFILLER_17_343 VPWR VGND sg13g2_fill_1
XFILLER_17_376 VPWR VGND sg13g2_decap_8
XFILLER_44_184 VPWR VGND sg13g2_fill_2
XFILLER_32_357 VPWR VGND sg13g2_fill_1
XFILLER_41_891 VPWR VGND sg13g2_decap_8
X_2710_ _0042_ _0966_ _0967_ VPWR VGND sg13g2_nand2_1
XFILLER_40_390 VPWR VGND sg13g2_fill_2
X_3690_ VGND VPWR net785 _0543_ _1660_ net770 sg13g2_a21oi_1
X_2641_ _0056_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[1\]
+ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\] _0912_ VPWR VGND sg13g2_nor4_1
X_2572_ _0858_ VPWR _0013_ VGND net583 _0857_ sg13g2_o21ai_1
XFILLER_5_792 VPWR VGND sg13g2_decap_8
X_4311_ net734 VGND VPWR net938 u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] clknet_leaf_47_clk
+ sg13g2_dfrbpq_2
X_4242_ net640 VGND VPWR net496 net31 clknet_leaf_0_clk sg13g2_dfrbpq_1
X_4173_ net660 VGND VPWR net217 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[9\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3124_ net329 net605 _1218_ VPWR VGND sg13g2_nor2_1
XFILLER_49_991 VPWR VGND sg13g2_decap_8
X_3055_ VGND VPWR net612 _1180_ _0189_ _1179_ sg13g2_a21oi_1
Xclkbuf_leaf_47_clk clknet_3_4__leaf_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
XFILLER_36_641 VPWR VGND sg13g2_fill_1
XFILLER_36_696 VPWR VGND sg13g2_decap_8
XFILLER_35_184 VPWR VGND sg13g2_fill_1
XFILLER_23_368 VPWR VGND sg13g2_fill_1
X_3957_ _1845_ _1846_ _1844_ _1847_ VPWR VGND sg13g2_nand3_1
X_2908_ net376 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ _1100_ _0122_ VPWR VGND sg13g2_mux2_1
X_3888_ _1961_ net382 net703 _1798_ VPWR VGND sg13g2_nor3_2
X_2839_ _1063_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] _1040_
+ VPWR VGND sg13g2_xnor2_1
Xfanout576 net577 net576 VPWR VGND sg13g2_buf_1
Xfanout587 net588 net587 VPWR VGND sg13g2_buf_2
Xfanout598 _0592_ net598 VPWR VGND sg13g2_buf_8
XFILLER_46_449 VPWR VGND sg13g2_fill_2
XFILLER_18_118 VPWR VGND sg13g2_decap_8
XFILLER_18_129 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_38_clk clknet_3_5__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_41_198 VPWR VGND sg13g2_fill_1
XFILLER_2_795 VPWR VGND sg13g2_decap_8
XFILLER_38_928 VPWR VGND sg13g2_decap_8
XFILLER_49_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_3_7__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_17_173 VPWR VGND sg13g2_fill_2
XFILLER_33_622 VPWR VGND sg13g2_fill_1
XFILLER_45_493 VPWR VGND sg13g2_decap_4
XFILLER_33_633 VPWR VGND sg13g2_fill_2
XFILLER_33_644 VPWR VGND sg13g2_fill_1
X_3811_ VGND VPWR net740 net318 _1744_ net331 sg13g2_a21oi_1
X_3742_ net763 net933 net589 _0365_ VPWR VGND sg13g2_mux2_1
X_3673_ _1643_ VPWR _1644_ VGND net992 net625 sg13g2_o21ai_1
X_2624_ _0024_ _0901_ _1956_ _0603_ _0592_ VPWR VGND sg13g2_a22oi_1
X_2555_ VGND VPWR _0844_ net585 _0626_ sg13g2_or2_1
X_2486_ _0676_ net617 _0747_ _0749_ _0783_ VPWR VGND sg13g2_nor4_1
X_4225_ net663 VGND VPWR net168 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[61\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
X_4156_ net672 VGND VPWR net998 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[0\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_2
X_3107_ _1209_ net197 _1202_ VPWR VGND sg13g2_nand2_1
X_4087_ net670 VGND VPWR net439 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[7\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_37_961 VPWR VGND sg13g2_decap_8
XFILLER_43_419 VPWR VGND sg13g2_fill_1
X_3038_ net546 net611 _1169_ VPWR VGND sg13g2_nor2_1
XFILLER_36_460 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_fill_2
XFILLER_24_677 VPWR VGND sg13g2_decap_8
XFILLER_24_688 VPWR VGND sg13g2_fill_2
XFILLER_11_327 VPWR VGND sg13g2_fill_2
XFILLER_11_65 VPWR VGND sg13g2_decap_4
XFILLER_19_427 VPWR VGND sg13g2_fill_2
XFILLER_47_758 VPWR VGND sg13g2_decap_8
XFILLER_46_235 VPWR VGND sg13g2_decap_8
XFILLER_43_964 VPWR VGND sg13g2_decap_8
XFILLER_7_810 VPWR VGND sg13g2_decap_8
X_2340_ _0641_ u_usb_cdc.u_ctrl_endp.state_q\[7\] _0640_ VPWR VGND sg13g2_nand2_1
XFILLER_2_592 VPWR VGND sg13g2_decap_8
X_2271_ _0573_ _1906_ _1986_ VPWR VGND sg13g2_nand2_2
XFILLER_42_1012 VPWR VGND sg13g2_decap_8
XFILLER_28_4 VPWR VGND sg13g2_fill_1
X_4010_ _1888_ net165 _1887_ VPWR VGND sg13g2_nand2_1
XFILLER_38_703 VPWR VGND sg13g2_decap_8
XFILLER_38_747 VPWR VGND sg13g2_fill_1
XFILLER_34_920 VPWR VGND sg13g2_fill_1
XFILLER_34_931 VPWR VGND sg13g2_decap_8
X_3725_ _1688_ VPWR _0351_ VGND _1899_ net598 sg13g2_o21ai_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_3656_ _1627_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[69\] net626
+ VPWR VGND sg13g2_nand2_1
X_3587_ net798 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[2\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[10\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[18\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[26\]
+ net791 _1561_ VPWR VGND sg13g2_mux4_1
X_2607_ _0888_ net762 u_usb_cdc.u_sie.data_q\[6\] VPWR VGND sg13g2_xnor2_1
X_2538_ _0008_ _0830_ _0831_ VPWR VGND sg13g2_nand2_1
XFILLER_0_507 VPWR VGND sg13g2_decap_8
X_4208_ net660 VGND VPWR net65 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[44\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_2469_ net720 net751 _0766_ VPWR VGND sg13g2_nor2_1
XFILLER_29_736 VPWR VGND sg13g2_fill_1
X_4139_ net650 VGND VPWR net494 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[59\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_44_717 VPWR VGND sg13g2_fill_1
XFILLER_43_205 VPWR VGND sg13g2_decap_4
XFILLER_16_419 VPWR VGND sg13g2_decap_4
XFILLER_37_791 VPWR VGND sg13g2_fill_1
XFILLER_24_441 VPWR VGND sg13g2_fill_2
XFILLER_24_452 VPWR VGND sg13g2_decap_8
XFILLER_40_956 VPWR VGND sg13g2_decap_8
XFILLER_12_669 VPWR VGND sg13g2_fill_2
XFILLER_7_139 VPWR VGND sg13g2_fill_1
XFILLER_4_802 VPWR VGND sg13g2_decap_8
XFILLER_4_879 VPWR VGND sg13g2_decap_8
XFILLER_47_522 VPWR VGND sg13g2_fill_2
XFILLER_19_268 VPWR VGND sg13g2_fill_2
XFILLER_19_279 VPWR VGND sg13g2_decap_8
XFILLER_35_728 VPWR VGND sg13g2_decap_4
XFILLER_15_474 VPWR VGND sg13g2_fill_1
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_31_989 VPWR VGND sg13g2_decap_8
X_3510_ _0338_ net573 _1486_ net576 _1938_ VPWR VGND sg13g2_a22oi_1
XFILLER_11_691 VPWR VGND sg13g2_fill_1
XFILLER_7_673 VPWR VGND sg13g2_decap_4
Xhold618 _0405_ VPWR VGND net936 sg13g2_dlygate4sd3_1
Xhold607 _0070_ VPWR VGND net925 sg13g2_dlygate4sd3_1
X_3441_ _1449_ net252 net580 VPWR VGND sg13g2_nand2_1
Xhold629 _0859_ VPWR VGND net947 sg13g2_dlygate4sd3_1
X_3372_ VGND VPWR net720 _1399_ _0285_ _1401_ sg13g2_a21oi_1
X_2323_ _0624_ _0610_ _0623_ VPWR VGND sg13g2_nand2_1
X_2254_ _0556_ _0049_ u_usb_cdc.u_ctrl_endp.state_q\[7\] VPWR VGND sg13g2_nand2b_1
X_2185_ _0486_ _0485_ u_usb_cdc.u_sie.data_q\[6\] _0487_ VPWR VGND sg13g2_mux2_1
XFILLER_25_205 VPWR VGND sg13g2_decap_8
XFILLER_26_706 VPWR VGND sg13g2_decap_8
XFILLER_21_455 VPWR VGND sg13g2_fill_2
XFILLER_22_989 VPWR VGND sg13g2_fill_2
X_3708_ _1676_ VPWR _1677_ VGND _1674_ _1675_ sg13g2_o21ai_1
X_3639_ _1610_ VPWR _1611_ VGND net799 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[36\]
+ sg13g2_o21ai_1
XFILLER_1_827 VPWR VGND sg13g2_decap_8
XFILLER_49_809 VPWR VGND sg13g2_decap_8
XFILLER_29_511 VPWR VGND sg13g2_fill_1
XFILLER_1_1009 VPWR VGND sg13g2_decap_8
XFILLER_44_558 VPWR VGND sg13g2_fill_1
XFILLER_40_720 VPWR VGND sg13g2_decap_8
XFILLER_13_978 VPWR VGND sg13g2_decap_8
XFILLER_9_938 VPWR VGND sg13g2_decap_8
XFILLER_33_74 VPWR VGND sg13g2_fill_2
XFILLER_4_676 VPWR VGND sg13g2_decap_8
XFILLER_39_308 VPWR VGND sg13g2_fill_2
XFILLER_0_871 VPWR VGND sg13g2_decap_8
Xhold4 u_usb_cdc.u_sie.u_phy_rx.dn_q\[1\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_48_875 VPWR VGND sg13g2_decap_8
XFILLER_16_761 VPWR VGND sg13g2_fill_1
X_3990_ net1001 VPWR _0431_ VGND _1825_ _1871_ sg13g2_o21ai_1
X_2941_ _1118_ net59 _1110_ VPWR VGND sg13g2_nand2_1
XFILLER_43_591 VPWR VGND sg13g2_fill_2
X_2872_ _1086_ net178 _1080_ VPWR VGND sg13g2_nand2_1
XFILLER_30_263 VPWR VGND sg13g2_fill_1
Xhold415 _0113_ VPWR VGND net457 sg13g2_dlygate4sd3_1
Xhold404 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[34\] VPWR VGND
+ net446 sg13g2_dlygate4sd3_1
Xhold426 _0119_ VPWR VGND net468 sg13g2_dlygate4sd3_1
Xhold437 u_usb_cdc.u_ctrl_endp.in_endp_q VPWR VGND net479 sg13g2_dlygate4sd3_1
Xhold459 _0220_ VPWR VGND net501 sg13g2_dlygate4sd3_1
X_3424_ _1439_ net772 _1424_ VPWR VGND sg13g2_nand2_1
Xhold448 _0108_ VPWR VGND net490 sg13g2_dlygate4sd3_1
X_3355_ net510 net570 _1392_ VPWR VGND sg13g2_nor2_1
X_3286_ _1351_ _1296_ net143 net602 net874 VPWR VGND sg13g2_a22oi_1
X_2306_ VGND VPWR _0607_ net749 u_usb_cdc.u_sie.out_eop_q sg13g2_or2_1
X_2237_ _0532_ _0533_ _0535_ _0539_ VPWR VGND sg13g2_nor3_1
X_2168_ net754 net758 _0470_ VPWR VGND sg13g2_xor2_1
X_2099_ VPWR _1977_ net466 VGND sg13g2_inv_1
XFILLER_41_539 VPWR VGND sg13g2_decap_4
XFILLER_10_904 VPWR VGND sg13g2_decap_8
XFILLER_6_919 VPWR VGND sg13g2_decap_8
XFILLER_1_624 VPWR VGND sg13g2_decap_8
XFILLER_29_330 VPWR VGND sg13g2_fill_1
XFILLER_28_63 VPWR VGND sg13g2_fill_1
XFILLER_45_856 VPWR VGND sg13g2_decap_8
XFILLER_17_558 VPWR VGND sg13g2_decap_4
XFILLER_44_95 VPWR VGND sg13g2_fill_1
XFILLER_5_974 VPWR VGND sg13g2_decap_8
XFILLER_4_451 VPWR VGND sg13g2_decap_8
X_3140_ _1226_ VPWR _0228_ VGND _1898_ net628 sg13g2_o21ai_1
X_3071_ _1190_ net204 net608 VPWR VGND sg13g2_nand2_1
X_2022_ _1901_ net752 VPWR VGND sg13g2_inv_8
XFILLER_36_889 VPWR VGND sg13g2_fill_2
X_3973_ _1861_ _1860_ _1806_ _1818_ net368 VPWR VGND sg13g2_a22oi_1
X_2924_ _1109_ net80 _1101_ VPWR VGND sg13g2_nand2_1
X_2855_ _1074_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net636 VPWR VGND sg13g2_nand2_1
XFILLER_8_790 VPWR VGND sg13g2_decap_4
Xhold201 _0199_ VPWR VGND net243 sg13g2_dlygate4sd3_1
X_2786_ u_usb_cdc.addr\[0\] _0870_ _1029_ VPWR VGND sg13g2_nor2_1
Xhold212 _0096_ VPWR VGND net254 sg13g2_dlygate4sd3_1
Xhold223 u_usb_cdc.u_sie.u_phy_tx.data_q\[3\] VPWR VGND net265 sg13g2_dlygate4sd3_1
Xhold234 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[50\] VPWR
+ VGND net276 sg13g2_dlygate4sd3_1
XFILLER_49_18 VPWR VGND sg13g2_decap_8
Xhold278 _0320_ VPWR VGND net320 sg13g2_dlygate4sd3_1
Xhold256 _0395_ VPWR VGND net298 sg13g2_dlygate4sd3_1
Xhold245 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[5\] VPWR VGND net287 sg13g2_dlygate4sd3_1
X_4456_ u_usb_cdc.out_valid_o[0] net22 VPWR VGND sg13g2_buf_1
Xhold267 _0073_ VPWR VGND net309 sg13g2_dlygate4sd3_1
Xhold289 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[1\] VPWR VGND net331 sg13g2_dlygate4sd3_1
X_4387_ net723 VGND VPWR net403 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[8\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xfanout703 _0449_ net703 VPWR VGND sg13g2_buf_8
Xfanout714 _1929_ net714 VPWR VGND sg13g2_buf_8
X_3407_ _1915_ _1424_ _1427_ VPWR VGND sg13g2_nor2_1
X_3338_ _1385_ net269 _1384_ VPWR VGND sg13g2_nand2_1
Xfanout758 net759 net758 VPWR VGND sg13g2_buf_8
Xfanout725 net727 net725 VPWR VGND sg13g2_buf_8
Xfanout747 net944 net747 VPWR VGND sg13g2_buf_8
Xfanout736 net737 net736 VPWR VGND sg13g2_buf_8
Xfanout769 net1056 net769 VPWR VGND sg13g2_buf_8
X_3269_ net329 net128 net814 _1335_ VPWR VGND sg13g2_mux2_1
XFILLER_39_672 VPWR VGND sg13g2_fill_1
XFILLER_14_517 VPWR VGND sg13g2_fill_1
XFILLER_41_325 VPWR VGND sg13g2_decap_4
XFILLER_6_716 VPWR VGND sg13g2_decap_8
XFILLER_2_900 VPWR VGND sg13g2_decap_8
XFILLER_30_42 VPWR VGND sg13g2_fill_2
XFILLER_1_421 VPWR VGND sg13g2_decap_8
XFILLER_7_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_977 VPWR VGND sg13g2_decap_8
XFILLER_1_498 VPWR VGND sg13g2_decap_8
XFILLER_44_130 VPWR VGND sg13g2_fill_1
XFILLER_44_174 VPWR VGND sg13g2_decap_4
XFILLER_33_837 VPWR VGND sg13g2_decap_8
XFILLER_40_380 VPWR VGND sg13g2_fill_1
XFILLER_9_576 VPWR VGND sg13g2_decap_4
X_2640_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[2\] u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[6\]
+ _0911_ VPWR VGND sg13g2_nor2_1
X_2571_ _0858_ _0646_ net871 _0638_ net866 VPWR VGND sg13g2_a22oi_1
XFILLER_5_771 VPWR VGND sg13g2_decap_8
X_4310_ net680 VGND VPWR net251 u_usb_cdc.u_sie.addr_q\[6\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_45_1010 VPWR VGND sg13g2_decap_8
X_4241_ net640 VGND VPWR net895 net30 clknet_leaf_55_clk sg13g2_dfrbpq_1
X_4172_ net660 VGND VPWR net105 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[8\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
XFILLER_49_970 VPWR VGND sg13g2_decap_8
X_3123_ VGND VPWR _1178_ net605 _0220_ net500 sg13g2_a21oi_1
X_3054_ _1180_ net752 net630 VPWR VGND sg13g2_nand2_2
XFILLER_36_631 VPWR VGND sg13g2_fill_2
XFILLER_11_509 VPWR VGND sg13g2_decap_8
XFILLER_23_358 VPWR VGND sg13g2_fill_2
X_3956_ _1846_ _1942_ u_usb_cdc.u_sie.phy_state_q\[4\] _1922_ net830 VPWR VGND sg13g2_a22oi_1
X_2907_ net475 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ _1100_ _0121_ VPWR VGND sg13g2_mux2_1
XFILLER_31_380 VPWR VGND sg13g2_decap_8
X_3887_ VGND VPWR net741 net264 _0404_ _1797_ sg13g2_a21oi_1
X_2838_ _1062_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2769_ net836 _0598_ _1004_ _1007_ _1014_ VPWR VGND sg13g2_and4_1
X_4439_ net698 VGND VPWR net313 _0059_ clknet_leaf_30_clk sg13g2_dfrbpq_1
Xfanout588 _0627_ net588 VPWR VGND sg13g2_buf_1
Xfanout599 _0972_ net599 VPWR VGND sg13g2_buf_8
Xfanout577 _1483_ net577 VPWR VGND sg13g2_buf_8
XFILLER_27_631 VPWR VGND sg13g2_fill_1
XFILLER_27_642 VPWR VGND sg13g2_fill_1
XFILLER_27_686 VPWR VGND sg13g2_decap_4
XFILLER_41_133 VPWR VGND sg13g2_fill_2
XFILLER_25_75 VPWR VGND sg13g2_decap_4
XFILLER_25_97 VPWR VGND sg13g2_fill_2
XFILLER_2_774 VPWR VGND sg13g2_decap_8
XFILLER_46_984 VPWR VGND sg13g2_decap_8
XFILLER_18_675 VPWR VGND sg13g2_fill_2
XFILLER_33_601 VPWR VGND sg13g2_fill_1
X_3810_ net712 _1742_ _1743_ VPWR VGND sg13g2_nor2_1
XFILLER_32_133 VPWR VGND sg13g2_fill_1
X_3741_ u_usb_cdc.u_sie.data_q\[1\] net962 net589 _0364_ VPWR VGND sg13g2_mux2_1
X_3672_ _1642_ VPWR _1643_ VGND _1529_ _1641_ sg13g2_o21ai_1
X_2623_ _0592_ VPWR _0901_ VGND net832 _0900_ sg13g2_o21ai_1
X_2554_ _0842_ VPWR _0001_ VGND _0741_ _0843_ sg13g2_o21ai_1
X_2485_ _0676_ _0747_ _0782_ VPWR VGND sg13g2_nor2_1
X_4224_ net664 VGND VPWR net249 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[60\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_1
X_4155_ net648 VGND VPWR _0158_ u_usb_cdc.in_ready_o[0] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3106_ _1208_ VPWR _0212_ VGND net709 _1161_ sg13g2_o21ai_1
XFILLER_28_417 VPWR VGND sg13g2_decap_8
X_4086_ net670 VGND VPWR net381 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[6\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_37_940 VPWR VGND sg13g2_decap_8
X_3037_ VGND VPWR net611 _1168_ _0183_ _1167_ sg13g2_a21oi_1
XFILLER_24_634 VPWR VGND sg13g2_decap_8
XFILLER_12_829 VPWR VGND sg13g2_fill_1
X_3939_ _1831_ _1828_ _1829_ _1830_ VPWR VGND sg13g2_and3_1
XFILLER_20_862 VPWR VGND sg13g2_fill_2
XFILLER_47_737 VPWR VGND sg13g2_decap_8
XFILLER_28_984 VPWR VGND sg13g2_decap_8
XFILLER_43_943 VPWR VGND sg13g2_decap_8
XFILLER_14_100 VPWR VGND sg13g2_fill_2
XFILLER_14_188 VPWR VGND sg13g2_fill_1
XFILLER_35_1020 VPWR VGND sg13g2_decap_8
XFILLER_10_350 VPWR VGND sg13g2_decap_8
XFILLER_7_899 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_8
XFILLER_2_571 VPWR VGND sg13g2_decap_8
X_2270_ _1906_ net706 _0572_ VPWR VGND sg13g2_and2_1
XFILLER_37_203 VPWR VGND sg13g2_decap_4
XFILLER_25_409 VPWR VGND sg13g2_decap_4
XFILLER_46_781 VPWR VGND sg13g2_decap_8
XFILLER_34_987 VPWR VGND sg13g2_decap_8
XFILLER_21_626 VPWR VGND sg13g2_decap_8
XFILLER_21_637 VPWR VGND sg13g2_fill_2
XFILLER_21_648 VPWR VGND sg13g2_fill_2
X_3724_ net590 _1683_ net980 _1688_ VPWR VGND sg13g2_nand3_1
X_3655_ _1626_ net995 net593 VPWR VGND sg13g2_nand2_1
X_2606_ _0887_ u_usb_cdc.u_sie.data_q\[3\] u_usb_cdc.u_sie.data_q\[7\] VPWR VGND sg13g2_xnor2_1
X_3586_ _1560_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[66\] net626
+ VPWR VGND sg13g2_nand2_1
X_2537_ net860 _0737_ _0799_ _0801_ _0831_ VPWR VGND sg13g2_or4_1
X_2468_ _0704_ _0705_ _0653_ _0765_ VPWR VGND sg13g2_nand3_1
X_4207_ net644 VGND VPWR net196 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[43\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2399_ _0699_ _0675_ net574 VPWR VGND sg13g2_nand2_1
XFILLER_29_726 VPWR VGND sg13g2_fill_1
X_4138_ net650 VGND VPWR net512 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[58\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_4069_ net691 VGND VPWR net220 u_usb_cdc.u_sie.addr_q\[0\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_25_965 VPWR VGND sg13g2_decap_4
XFILLER_40_935 VPWR VGND sg13g2_decap_8
XFILLER_11_114 VPWR VGND sg13g2_decap_4
XFILLER_25_998 VPWR VGND sg13g2_decap_8
XFILLER_11_125 VPWR VGND sg13g2_fill_1
XFILLER_11_136 VPWR VGND sg13g2_decap_8
XFILLER_7_129 VPWR VGND sg13g2_fill_1
XFILLER_22_87 VPWR VGND sg13g2_fill_1
XFILLER_4_858 VPWR VGND sg13g2_decap_8
XFILLER_3_313 VPWR VGND sg13g2_fill_2
XFILLER_26_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_501 VPWR VGND sg13g2_decap_8
XFILLER_47_589 VPWR VGND sg13g2_fill_1
XFILLER_19_258 VPWR VGND sg13g2_fill_1
XFILLER_31_968 VPWR VGND sg13g2_decap_8
XFILLER_10_180 VPWR VGND sg13g2_fill_1
Xhold608 u_usb_cdc.addr\[2\] VPWR VGND net926 sg13g2_dlygate4sd3_1
Xhold619 u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] VPWR VGND net937 sg13g2_dlygate4sd3_1
X_3440_ VGND VPWR _1908_ _0869_ _0306_ _1448_ sg13g2_a21oi_1
X_3371_ net910 _1399_ _1401_ VPWR VGND sg13g2_nor2_1
XFILLER_40_4 VPWR VGND sg13g2_decap_4
X_2322_ _1924_ _0468_ _0623_ VPWR VGND sg13g2_nor2_2
X_2253_ u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\] u_usb_cdc.u_ctrl_endp.req_q\[4\] _0555_
+ VPWR VGND sg13g2_nor2b_1
X_2184_ _0472_ u_usb_cdc.u_sie.data_q\[4\] _0486_ VPWR VGND sg13g2_xor2_1
XFILLER_22_902 VPWR VGND sg13g2_decap_8
XFILLER_34_740 VPWR VGND sg13g2_fill_1
XFILLER_33_261 VPWR VGND sg13g2_fill_2
XFILLER_34_773 VPWR VGND sg13g2_fill_2
XFILLER_22_979 VPWR VGND sg13g2_fill_2
XFILLER_21_467 VPWR VGND sg13g2_decap_4
X_3707_ VGND VPWR _1668_ _1670_ _1676_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\]
+ sg13g2_a21oi_1
XFILLER_49_1019 VPWR VGND sg13g2_decap_8
X_3638_ VGND VPWR net799 _1971_ _1610_ net793 sg13g2_a21oi_1
XFILLER_1_806 VPWR VGND sg13g2_decap_8
X_3569_ VGND VPWR _1544_ _0705_ net776 sg13g2_or2_1
XFILLER_29_545 VPWR VGND sg13g2_fill_2
XFILLER_29_567 VPWR VGND sg13g2_fill_2
XFILLER_24_250 VPWR VGND sg13g2_fill_2
XFILLER_40_743 VPWR VGND sg13g2_fill_1
XFILLER_9_917 VPWR VGND sg13g2_decap_8
XFILLER_13_957 VPWR VGND sg13g2_decap_8
XFILLER_12_456 VPWR VGND sg13g2_decap_4
XFILLER_4_611 VPWR VGND sg13g2_decap_8
XFILLER_4_655 VPWR VGND sg13g2_decap_8
XFILLER_3_132 VPWR VGND sg13g2_decap_4
XFILLER_0_850 VPWR VGND sg13g2_decap_8
XFILLER_48_854 VPWR VGND sg13g2_decap_8
Xhold5 u_usb_cdc.u_sie.u_phy_rx.dp_q\[1\] VPWR VGND net47 sg13g2_dlygate4sd3_1
X_2940_ _1117_ VPWR _0137_ VGND _1965_ _1095_ sg13g2_o21ai_1
XFILLER_43_570 VPWR VGND sg13g2_decap_8
XFILLER_16_784 VPWR VGND sg13g2_decap_4
XFILLER_31_732 VPWR VGND sg13g2_fill_2
X_2871_ _1084_ VPWR _0100_ VGND net826 _1085_ sg13g2_o21ai_1
Xhold405 _0117_ VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold416 u_usb_cdc.u_ctrl_endp.addr_dd\[5\] VPWR VGND net458 sg13g2_dlygate4sd3_1
XFILLER_8_994 VPWR VGND sg13g2_decap_8
Xhold427 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[70\] VPWR VGND
+ net469 sg13g2_dlygate4sd3_1
Xhold438 _0267_ VPWR VGND net480 sg13g2_dlygate4sd3_1
X_3423_ _1436_ VPWR _0299_ VGND _1426_ _1438_ sg13g2_o21ai_1
Xhold449 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[71\] VPWR VGND
+ net491 sg13g2_dlygate4sd3_1
X_3354_ VGND VPWR net718 net571 _0277_ _1391_ sg13g2_a21oi_1
X_3285_ net805 net602 _1349_ _1350_ VPWR VGND sg13g2_nor3_1
X_2305_ net749 _0605_ _0606_ VPWR VGND sg13g2_nor2_2
X_2236_ net787 u_usb_cdc.u_ctrl_endp.max_length_q\[0\] _0538_ VPWR VGND sg13g2_xor2_1
XFILLER_39_854 VPWR VGND sg13g2_fill_1
X_2167_ net1009 _0466_ _0468_ _0469_ VPWR VGND sg13g2_or3_1
X_2098_ VPWR _1976_ net265 VGND sg13g2_inv_1
XFILLER_21_264 VPWR VGND sg13g2_fill_2
XFILLER_1_603 VPWR VGND sg13g2_decap_8
XFILLER_29_364 VPWR VGND sg13g2_decap_4
XFILLER_45_835 VPWR VGND sg13g2_decap_8
XFILLER_44_301 VPWR VGND sg13g2_fill_1
XFILLER_44_345 VPWR VGND sg13g2_fill_2
XFILLER_32_518 VPWR VGND sg13g2_decap_4
XFILLER_9_714 VPWR VGND sg13g2_decap_4
XFILLER_9_769 VPWR VGND sg13g2_fill_1
XFILLER_40_584 VPWR VGND sg13g2_fill_2
XFILLER_5_953 VPWR VGND sg13g2_decap_8
XFILLER_5_79 VPWR VGND sg13g2_decap_8
X_3070_ _1189_ VPWR _0195_ VGND _1899_ net609 sg13g2_o21ai_1
XFILLER_48_662 VPWR VGND sg13g2_decap_4
X_2021_ net751 _1900_ VPWR VGND sg13g2_inv_4
XFILLER_48_695 VPWR VGND sg13g2_fill_2
XFILLER_47_161 VPWR VGND sg13g2_fill_2
XFILLER_36_879 VPWR VGND sg13g2_fill_1
XFILLER_35_389 VPWR VGND sg13g2_decap_4
XFILLER_16_592 VPWR VGND sg13g2_decap_8
X_3972_ VGND VPWR _1808_ _1859_ _1860_ _1818_ sg13g2_a21oi_1
X_2923_ _1108_ VPWR _0129_ VGND _1076_ _1099_ sg13g2_o21ai_1
X_2854_ _1073_ net253 _1059_ VPWR VGND sg13g2_nand2_1
X_2785_ _0071_ _1028_ _1023_ _1026_ net355 VPWR VGND sg13g2_a22oi_1
Xhold202 u_usb_cdc.u_sie.u_phy_rx.se0_q VPWR VGND net244 sg13g2_dlygate4sd3_1
Xhold224 _0424_ VPWR VGND net266 sg13g2_dlygate4sd3_1
Xhold213 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[0\] VPWR VGND
+ net255 sg13g2_dlygate4sd3_1
Xhold235 _0217_ VPWR VGND net277 sg13g2_dlygate4sd3_1
Xhold257 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[20\] VPWR
+ VGND net299 sg13g2_dlygate4sd3_1
Xhold246 _0386_ VPWR VGND net288 sg13g2_dlygate4sd3_1
Xhold268 u_usb_cdc.u_sie.in_toggle_q\[0\] VPWR VGND net310 sg13g2_dlygate4sd3_1
Xhold279 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[18\] VPWR
+ VGND net321 sg13g2_dlygate4sd3_1
X_4386_ net723 VGND VPWR _0388_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[7\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xfanout704 _0449_ net704 VPWR VGND sg13g2_buf_2
Xfanout715 _1916_ net715 VPWR VGND sg13g2_buf_8
X_3406_ _0844_ _1424_ _1425_ _1426_ VPWR VGND sg13g2_or3_1
Xfanout726 net733 net726 VPWR VGND sg13g2_buf_8
X_3337_ _0614_ _0639_ _1383_ _1384_ VPWR VGND sg13g2_nor3_2
Xfanout737 u_usb_cdc.clk_gate_q net737 VPWR VGND sg13g2_buf_8
Xfanout748 net944 net748 VPWR VGND sg13g2_buf_2
Xfanout759 u_usb_cdc.sie_out_data\[1\] net759 VPWR VGND sg13g2_buf_8
X_3268_ _1333_ VPWR _1334_ VGND net814 net139 sg13g2_o21ai_1
X_2219_ _0511_ _0505_ _0521_ VPWR VGND sg13g2_xor2_1
X_3199_ _1272_ _0606_ _1271_ net960 net749 VPWR VGND sg13g2_a22oi_1
XFILLER_38_194 VPWR VGND sg13g2_fill_2
XFILLER_5_205 VPWR VGND sg13g2_decap_4
XFILLER_30_54 VPWR VGND sg13g2_decap_8
XFILLER_30_65 VPWR VGND sg13g2_fill_1
XFILLER_1_400 VPWR VGND sg13g2_decap_8
XFILLER_2_956 VPWR VGND sg13g2_decap_8
XFILLER_1_477 VPWR VGND sg13g2_decap_8
XFILLER_18_846 VPWR VGND sg13g2_decap_8
XFILLER_45_687 VPWR VGND sg13g2_decap_8
XFILLER_44_142 VPWR VGND sg13g2_fill_1
XFILLER_26_890 VPWR VGND sg13g2_fill_1
XFILLER_13_573 VPWR VGND sg13g2_decap_8
XFILLER_40_392 VPWR VGND sg13g2_fill_1
XFILLER_5_750 VPWR VGND sg13g2_decap_8
X_2570_ _0857_ net550 _0856_ VPWR VGND sg13g2_nand2_1
X_4240_ net640 VGND VPWR net406 net29 clknet_leaf_1_clk sg13g2_dfrbpq_1
X_4171_ net662 VGND VPWR _0174_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[7\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3122_ net499 _1211_ _1217_ VPWR VGND sg13g2_nor2_1
X_3053_ net267 net612 _1179_ VPWR VGND sg13g2_nor2_1
XFILLER_36_665 VPWR VGND sg13g2_fill_2
X_3955_ _1845_ _1948_ net831 u_usb_cdc.u_sie.data_q\[4\] net834 VPWR VGND sg13g2_a22oi_1
X_2906_ net513 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ _1100_ _0120_ VPWR VGND sg13g2_mux2_1
X_3886_ net748 net741 _1797_ VPWR VGND sg13g2_nor2_1
X_2837_ net827 net828 _1061_ VPWR VGND sg13g2_nor2b_2
X_2768_ _0598_ _1004_ net836 _1013_ VPWR VGND _1007_ sg13g2_nand4_1
X_2699_ _0959_ net970 _0832_ VPWR VGND sg13g2_nand2_1
X_4438_ net698 VGND VPWR _0429_ _0058_ clknet_leaf_29_clk sg13g2_dfrbpq_2
X_4369_ net692 VGND VPWR net293 u_usb_cdc.u_sie.out_eop_q clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_47_919 VPWR VGND sg13g2_decap_8
Xfanout567 net568 net567 VPWR VGND sg13g2_buf_8
Xfanout589 _0602_ net589 VPWR VGND sg13g2_buf_8
Xfanout578 _1254_ net578 VPWR VGND sg13g2_buf_8
XFILLER_27_654 VPWR VGND sg13g2_fill_1
XFILLER_15_827 VPWR VGND sg13g2_fill_1
XFILLER_26_153 VPWR VGND sg13g2_decap_8
XFILLER_15_849 VPWR VGND sg13g2_fill_2
XFILLER_10_532 VPWR VGND sg13g2_decap_4
XFILLER_10_554 VPWR VGND sg13g2_fill_2
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_753 VPWR VGND sg13g2_decap_8
XFILLER_1_274 VPWR VGND sg13g2_decap_8
XFILLER_37_418 VPWR VGND sg13g2_fill_2
XFILLER_37_407 VPWR VGND sg13g2_fill_2
XFILLER_46_963 VPWR VGND sg13g2_decap_8
XFILLER_17_153 VPWR VGND sg13g2_fill_1
XFILLER_18_665 VPWR VGND sg13g2_decap_4
XFILLER_13_370 VPWR VGND sg13g2_decap_8
XFILLER_14_882 VPWR VGND sg13g2_decap_8
XFILLER_20_307 VPWR VGND sg13g2_fill_1
X_3740_ u_usb_cdc.u_sie.data_q\[0\] net911 net589 _0363_ VPWR VGND sg13g2_mux2_1
XFILLER_32_178 VPWR VGND sg13g2_decap_4
XFILLER_12_1021 VPWR VGND sg13g2_decap_4
X_3671_ VGND VPWR net631 _1635_ _1642_ _1489_ sg13g2_a21oi_1
X_2622_ _0891_ _0899_ _0900_ VPWR VGND sg13g2_nor2_1
X_2553_ _0843_ _0795_ _0794_ VPWR VGND sg13g2_nand2b_1
X_2484_ _1933_ _0686_ _0713_ _0743_ _0781_ VPWR VGND sg13g2_nor4_1
X_4223_ net644 VGND VPWR _0226_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[59\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_4154_ net683 VGND VPWR net902 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_29_908 VPWR VGND sg13g2_decap_4
X_4085_ net651 VGND VPWR net555 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[5\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3105_ _1208_ net108 _1202_ VPWR VGND sg13g2_nand2_1
X_3036_ _1168_ net761 net630 VPWR VGND sg13g2_nand2_2
XFILLER_36_440 VPWR VGND sg13g2_fill_1
XFILLER_37_996 VPWR VGND sg13g2_decap_8
XFILLER_11_329 VPWR VGND sg13g2_fill_1
XFILLER_23_167 VPWR VGND sg13g2_fill_1
X_3938_ _1830_ _1950_ net831 _1940_ net838 VPWR VGND sg13g2_a22oi_1
X_3869_ VGND VPWR _1784_ _1786_ _0397_ _1785_ sg13g2_a21oi_1
XFILLER_47_716 VPWR VGND sg13g2_decap_8
XFILLER_4_1019 VPWR VGND sg13g2_decap_4
XFILLER_28_963 VPWR VGND sg13g2_decap_8
XFILLER_43_922 VPWR VGND sg13g2_decap_8
XFILLER_15_624 VPWR VGND sg13g2_fill_1
XFILLER_27_495 VPWR VGND sg13g2_decap_8
XFILLER_43_999 VPWR VGND sg13g2_decap_8
XFILLER_42_476 VPWR VGND sg13g2_fill_2
XFILLER_10_340 VPWR VGND sg13g2_fill_1
XFILLER_7_878 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_37_237 VPWR VGND sg13g2_fill_2
XFILLER_46_760 VPWR VGND sg13g2_decap_8
XFILLER_34_966 VPWR VGND sg13g2_decap_8
X_3723_ _1687_ VPWR _0350_ VGND _1896_ net598 sg13g2_o21ai_1
XFILLER_20_159 VPWR VGND sg13g2_fill_2
X_3654_ _1604_ VPWR _0343_ VGND _1624_ _1625_ sg13g2_o21ai_1
X_2605_ _0886_ net764 u_usb_cdc.u_sie.data_q\[5\] VPWR VGND sg13g2_xnor2_1
X_3585_ _1559_ net763 net594 VPWR VGND sg13g2_nand2_1
X_2536_ net921 VPWR _0830_ VGND _0820_ _0829_ sg13g2_o21ai_1
X_2467_ _0688_ _0763_ u_usb_cdc.u_ctrl_endp.req_q\[6\] _0764_ VPWR VGND sg13g2_nand3_1
X_4206_ net645 VGND VPWR net133 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[42\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_2398_ net587 net584 net619 _0698_ VGND VPWR _0697_ sg13g2_nor4_2
X_4137_ net648 VGND VPWR net435 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[57\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_4068_ net699 VGND VPWR _0038_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
X_3019_ _1156_ net102 _1146_ VPWR VGND sg13g2_nand2_1
XFILLER_25_933 VPWR VGND sg13g2_fill_1
XFILLER_19_1016 VPWR VGND sg13g2_decap_8
XFILLER_19_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_914 VPWR VGND sg13g2_decap_8
XFILLER_12_649 VPWR VGND sg13g2_fill_2
XFILLER_4_837 VPWR VGND sg13g2_decap_8
XFILLER_47_524 VPWR VGND sg13g2_fill_1
XFILLER_47_557 VPWR VGND sg13g2_decap_8
XFILLER_27_270 VPWR VGND sg13g2_fill_1
XFILLER_42_251 VPWR VGND sg13g2_fill_2
XFILLER_15_465 VPWR VGND sg13g2_decap_8
XFILLER_30_424 VPWR VGND sg13g2_decap_8
XFILLER_30_468 VPWR VGND sg13g2_fill_1
Xhold609 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[1\] VPWR VGND
+ net927 sg13g2_dlygate4sd3_1
X_3370_ VGND VPWR net721 _1399_ _0284_ _1400_ sg13g2_a21oi_1
XFILLER_3_892 VPWR VGND sg13g2_decap_8
X_2321_ VGND VPWR _0620_ _0621_ _0622_ _0573_ sg13g2_a21oi_1
X_2252_ VPWR VGND _0553_ _0546_ _0551_ _0539_ _0554_ _0540_ sg13g2_a221oi_1
XFILLER_33_4 VPWR VGND sg13g2_decap_8
X_2183_ _0485_ _0483_ _0484_ VPWR VGND sg13g2_xnor2_1
XFILLER_46_590 VPWR VGND sg13g2_fill_1
XFILLER_22_914 VPWR VGND sg13g2_decap_8
XFILLER_33_273 VPWR VGND sg13g2_decap_8
X_3706_ net789 VPWR _1675_ VGND net793 _1672_ sg13g2_o21ai_1
XFILLER_30_991 VPWR VGND sg13g2_decap_8
X_3637_ _1608_ VPWR _1609_ VGND net793 _1606_ sg13g2_o21ai_1
X_3568_ net778 VPWR _1543_ VGND _0705_ _1542_ sg13g2_o21ai_1
X_2519_ _0815_ _0813_ _0814_ VPWR VGND sg13g2_nand2_1
X_3499_ _0328_ net572 net549 net575 _1950_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_339 VPWR VGND sg13g2_decap_8
XFILLER_17_719 VPWR VGND sg13g2_decap_4
XFILLER_25_741 VPWR VGND sg13g2_fill_2
XFILLER_13_936 VPWR VGND sg13g2_decap_8
XFILLER_33_32 VPWR VGND sg13g2_decap_8
XFILLER_40_777 VPWR VGND sg13g2_decap_4
XFILLER_8_428 VPWR VGND sg13g2_fill_2
XFILLER_32_1013 VPWR VGND sg13g2_decap_8
XFILLER_33_76 VPWR VGND sg13g2_fill_1
XFILLER_4_623 VPWR VGND sg13g2_fill_1
XFILLER_48_833 VPWR VGND sg13g2_decap_8
Xhold6 u_usb_cdc.clk_cnt_q\[0\] VPWR VGND net48 sg13g2_dlygate4sd3_1
XFILLER_35_538 VPWR VGND sg13g2_fill_2
XFILLER_35_549 VPWR VGND sg13g2_fill_2
XFILLER_15_262 VPWR VGND sg13g2_decap_4
X_2870_ _1085_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ _1082_ VPWR VGND sg13g2_nand2_1
XFILLER_31_777 VPWR VGND sg13g2_decap_8
XFILLER_31_788 VPWR VGND sg13g2_fill_1
XFILLER_8_973 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_3_2__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
Xhold417 _0280_ VPWR VGND net459 sg13g2_dlygate4sd3_1
Xhold406 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[68\] VPWR VGND
+ net448 sg13g2_dlygate4sd3_1
X_3422_ _1434_ net775 _1438_ VPWR VGND sg13g2_xor2_1
Xhold428 _0153_ VPWR VGND net470 sg13g2_dlygate4sd3_1
Xhold439 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[28\] VPWR VGND
+ net481 sg13g2_dlygate4sd3_1
X_3353_ net392 net570 _1391_ VPWR VGND sg13g2_nor2_1
X_3284_ VPWR VGND _1279_ _1347_ _1348_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[2\]
+ _1349_ _1344_ sg13g2_a221oi_1
XFILLER_24_0 VPWR VGND sg13g2_fill_1
X_2304_ net747 _0604_ _0605_ VPWR VGND sg13g2_nor2_2
X_2235_ net784 u_usb_cdc.u_ctrl_endp.max_length_q\[2\] _0537_ VPWR VGND sg13g2_xor2_1
X_2166_ _0468_ net1018 _0467_ VPWR VGND sg13g2_nand2_1
XFILLER_39_866 VPWR VGND sg13g2_fill_2
XFILLER_0_1011 VPWR VGND sg13g2_decap_8
XFILLER_26_538 VPWR VGND sg13g2_fill_1
XFILLER_19_590 VPWR VGND sg13g2_decap_4
X_2097_ _1975_ net979 VPWR VGND sg13g2_inv_2
XFILLER_41_508 VPWR VGND sg13g2_decap_4
XFILLER_22_755 VPWR VGND sg13g2_decap_8
XFILLER_22_766 VPWR VGND sg13g2_fill_2
X_2999_ _1142_ VPWR _0171_ VGND _1899_ net613 sg13g2_o21ai_1
XFILLER_10_939 VPWR VGND sg13g2_decap_8
XFILLER_1_659 VPWR VGND sg13g2_decap_8
XFILLER_49_608 VPWR VGND sg13g2_decap_4
XFILLER_45_814 VPWR VGND sg13g2_decap_8
XFILLER_44_357 VPWR VGND sg13g2_decap_4
XFILLER_13_722 VPWR VGND sg13g2_fill_2
XFILLER_25_571 VPWR VGND sg13g2_decap_4
XFILLER_12_254 VPWR VGND sg13g2_fill_1
XFILLER_8_269 VPWR VGND sg13g2_decap_8
XFILLER_5_932 VPWR VGND sg13g2_decap_8
X_2020_ net754 _1899_ VPWR VGND sg13g2_inv_4
XFILLER_36_814 VPWR VGND sg13g2_fill_2
XFILLER_35_324 VPWR VGND sg13g2_decap_4
XFILLER_39_1008 VPWR VGND sg13g2_decap_8
X_3971_ _1857_ _1858_ _0895_ _1859_ VPWR VGND sg13g2_nand3_1
X_2922_ _1108_ net71 _1101_ VPWR VGND sg13g2_nand2_1
XFILLER_31_552 VPWR VGND sg13g2_decap_8
X_2853_ _1071_ VPWR _0095_ VGND net616 _1072_ sg13g2_o21ai_1
X_2784_ _1932_ VPWR _1028_ VGND u_usb_cdc.u_ctrl_endp.endp_q\[0\] _1027_ sg13g2_o21ai_1
Xhold214 _0167_ VPWR VGND net256 sg13g2_dlygate4sd3_1
Xhold225 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[22\] VPWR
+ VGND net267 sg13g2_dlygate4sd3_1
Xhold203 _0432_ VPWR VGND net245 sg13g2_dlygate4sd3_1
Xhold247 u_usb_cdc.u_sie.in_byte_q\[0\] VPWR VGND net289 sg13g2_dlygate4sd3_1
Xhold258 _0187_ VPWR VGND net300 sg13g2_dlygate4sd3_1
Xhold236 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[4\] VPWR VGND net278 sg13g2_dlygate4sd3_1
Xhold269 _0069_ VPWR VGND net311 sg13g2_dlygate4sd3_1
Xfanout705 _2002_ net705 VPWR VGND sg13g2_buf_8
X_4385_ net722 VGND VPWR net173 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[6\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_3405_ VGND VPWR _0558_ _0605_ _1425_ u_usb_cdc.u_ctrl_endp.state_q\[6\] sg13g2_a21oi_1
X_3336_ u_usb_cdc.u_ctrl_endp.req_q\[7\] net841 _1383_ VPWR VGND sg13g2_nor2b_1
Xfanout727 net733 net727 VPWR VGND sg13g2_buf_8
Xfanout738 net739 net738 VPWR VGND sg13g2_buf_8
Xfanout749 net1068 net749 VPWR VGND sg13g2_buf_8
Xfanout716 _1916_ net716 VPWR VGND sg13g2_buf_1
X_3267_ _1333_ net814 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[46\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_27_803 VPWR VGND sg13g2_fill_2
X_2218_ _0520_ _0500_ net541 VPWR VGND sg13g2_xnor2_1
X_3198_ _1270_ VPWR _1271_ VGND net768 _1964_ sg13g2_o21ai_1
X_2149_ _0443_ _0447_ _0451_ _0452_ VPWR VGND sg13g2_nor3_1
XFILLER_42_828 VPWR VGND sg13g2_fill_1
XFILLER_14_508 VPWR VGND sg13g2_decap_8
XFILLER_26_368 VPWR VGND sg13g2_decap_8
XFILLER_14_56 VPWR VGND sg13g2_fill_2
XFILLER_30_44 VPWR VGND sg13g2_fill_1
XFILLER_2_935 VPWR VGND sg13g2_decap_8
XFILLER_1_456 VPWR VGND sg13g2_decap_8
XFILLER_45_600 VPWR VGND sg13g2_fill_1
XFILLER_29_140 VPWR VGND sg13g2_decap_4
XFILLER_13_530 VPWR VGND sg13g2_decap_8
XFILLER_9_523 VPWR VGND sg13g2_decap_4
X_4170_ net644 VGND VPWR net55 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[6\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3121_ VGND VPWR _1176_ net605 _0219_ _1216_ sg13g2_a21oi_1
X_3052_ VGND VPWR net612 _1178_ _0188_ _1177_ sg13g2_a21oi_1
XFILLER_36_633 VPWR VGND sg13g2_fill_1
XFILLER_35_154 VPWR VGND sg13g2_decap_8
X_3954_ _1844_ _1990_ _0579_ VPWR VGND sg13g2_nand2_1
X_3885_ VGND VPWR net741 _0975_ _0403_ net358 sg13g2_a21oi_1
X_2905_ net467 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ _1100_ _0119_ VPWR VGND sg13g2_mux2_1
X_2836_ _1060_ net95 _1059_ VPWR VGND sg13g2_nand2_1
X_2767_ VGND VPWR _1966_ _1010_ _0069_ _1012_ sg13g2_a21oi_1
XFILLER_2_209 VPWR VGND sg13g2_fill_1
X_2698_ _0038_ _0957_ net562 VPWR VGND sg13g2_nand2_1
X_4437_ net696 VGND VPWR net369 _0057_ clknet_leaf_28_clk sg13g2_dfrbpq_1
X_4368_ net692 VGND VPWR _0370_ u_usb_cdc.sie_out_err clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3319_ VGND VPWR _1913_ _1358_ _0261_ _1372_ sg13g2_a21oi_1
Xfanout568 _1406_ net568 VPWR VGND sg13g2_buf_8
X_4299_ net668 VGND VPWR net952 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
Xfanout579 _0933_ net579 VPWR VGND sg13g2_buf_8
XFILLER_39_460 VPWR VGND sg13g2_fill_2
XFILLER_23_883 VPWR VGND sg13g2_fill_2
XFILLER_25_99 VPWR VGND sg13g2_fill_1
XFILLER_22_382 VPWR VGND sg13g2_decap_4
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_10_588 VPWR VGND sg13g2_fill_2
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_29_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_257 VPWR VGND sg13g2_decap_8
XFILLER_2_48 VPWR VGND sg13g2_fill_1
XFILLER_38_909 VPWR VGND sg13g2_fill_2
XFILLER_46_942 VPWR VGND sg13g2_decap_8
XFILLER_12_1000 VPWR VGND sg13g2_decap_8
X_3670_ _1641_ _1638_ _1640_ _1573_ u_usb_cdc.u_ctrl_endp.req_q\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_9_397 VPWR VGND sg13g2_fill_2
X_2621_ net837 VPWR _0899_ VGND net764 _0890_ sg13g2_o21ai_1
X_2552_ net552 VPWR _0842_ VGND _0840_ _0841_ sg13g2_o21ai_1
X_4222_ net659 VGND VPWR _0225_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[58\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_2483_ _1933_ _0686_ _0780_ VPWR VGND sg13g2_nor2_1
X_4153_ net683 VGND VPWR _0156_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[2\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3104_ _1207_ VPWR _0211_ VGND net708 _1159_ sg13g2_o21ai_1
X_4084_ net654 VGND VPWR net398 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[4\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3035_ net389 net611 _1167_ VPWR VGND sg13g2_nor2_1
XFILLER_37_975 VPWR VGND sg13g2_decap_8
XFILLER_36_474 VPWR VGND sg13g2_decap_8
XFILLER_23_146 VPWR VGND sg13g2_fill_2
X_3937_ _1829_ net762 net834 u_usb_cdc.u_sie.pid_q\[2\] net830 VPWR VGND sg13g2_a22oi_1
X_3868_ _1782_ net566 _1740_ _1786_ VPWR VGND sg13g2_a21o_1
XFILLER_20_897 VPWR VGND sg13g2_fill_1
X_2819_ net4 net1032 net637 _0077_ VPWR VGND sg13g2_mux2_1
X_3799_ _1734_ net360 net579 VPWR VGND sg13g2_nand2_1
XFILLER_46_249 VPWR VGND sg13g2_fill_1
XFILLER_43_901 VPWR VGND sg13g2_decap_8
XFILLER_43_978 VPWR VGND sg13g2_decap_8
XFILLER_14_135 VPWR VGND sg13g2_decap_8
XFILLER_15_658 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_fill_2
XFILLER_7_824 VPWR VGND sg13g2_decap_8
XFILLER_7_857 VPWR VGND sg13g2_decap_8
XFILLER_42_1026 VPWR VGND sg13g2_fill_2
XFILLER_38_717 VPWR VGND sg13g2_fill_2
XFILLER_18_452 VPWR VGND sg13g2_decap_8
XFILLER_19_964 VPWR VGND sg13g2_decap_8
XFILLER_18_496 VPWR VGND sg13g2_decap_8
XFILLER_34_945 VPWR VGND sg13g2_decap_8
X_3722_ net590 _1683_ net1011 _1687_ VPWR VGND sg13g2_nand3_1
X_3653_ net597 VPWR _1625_ VGND net929 net624 sg13g2_o21ai_1
X_2604_ _0885_ net766 u_usb_cdc.u_sie.data_q\[4\] VPWR VGND sg13g2_xnor2_1
X_3584_ net594 net765 _1558_ _0340_ VPWR VGND sg13g2_a21o_1
X_2535_ _0821_ _0828_ _0712_ _0829_ VPWR VGND sg13g2_nand3_1
X_2466_ u_usb_cdc.u_ctrl_endp.rec_q\[1\] net618 _1926_ _0763_ VPWR VGND sg13g2_nand3_1
X_4205_ net659 VGND VPWR net247 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[41\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_2397_ _0697_ net738 _0688_ VPWR VGND sg13g2_nand2_1
X_4136_ net649 VGND VPWR net396 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[56\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_28_238 VPWR VGND sg13g2_decap_4
X_4067_ net698 VGND VPWR net383 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
XFILLER_37_761 VPWR VGND sg13g2_decap_8
X_3018_ _1154_ VPWR _0177_ VGND net821 _1155_ sg13g2_o21ai_1
XFILLER_7_109 VPWR VGND sg13g2_decap_8
XFILLER_4_816 VPWR VGND sg13g2_decap_8
XFILLER_3_315 VPWR VGND sg13g2_fill_1
XFILLER_3_337 VPWR VGND sg13g2_decap_4
XFILLER_47_536 VPWR VGND sg13g2_decap_8
XFILLER_27_260 VPWR VGND sg13g2_fill_1
XFILLER_42_230 VPWR VGND sg13g2_decap_8
XFILLER_27_293 VPWR VGND sg13g2_decap_4
XFILLER_43_786 VPWR VGND sg13g2_fill_1
XFILLER_8_58 VPWR VGND sg13g2_fill_1
XFILLER_7_687 VPWR VGND sg13g2_fill_2
XFILLER_3_871 VPWR VGND sg13g2_decap_8
X_2320_ u_usb_cdc.sie_in_data_ack u_usb_cdc.sie_in_req _0621_ VPWR VGND sg13g2_nor2_2
XFILLER_2_392 VPWR VGND sg13g2_decap_8
X_2251_ _0553_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] u_usb_cdc.u_ctrl_endp.req_q\[8\]
+ _0552_ VPWR VGND sg13g2_and3_1
X_2182_ _0484_ net764 _0470_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_536 VPWR VGND sg13g2_decap_8
XFILLER_38_558 VPWR VGND sg13g2_decap_8
XFILLER_21_403 VPWR VGND sg13g2_decap_8
XFILLER_33_263 VPWR VGND sg13g2_fill_1
XFILLER_34_775 VPWR VGND sg13g2_fill_1
XFILLER_30_970 VPWR VGND sg13g2_decap_8
X_3705_ VGND VPWR net801 _1974_ _1674_ _1673_ sg13g2_a21oi_1
X_3636_ VGND VPWR net796 _1607_ _1608_ net790 sg13g2_a21oi_1
X_3567_ _0660_ net781 _1542_ VPWR VGND sg13g2_nor2b_1
X_2518_ net618 _0782_ _0695_ _0814_ VPWR VGND sg13g2_nand3_1
X_3498_ _0327_ net572 net445 net575 _1951_ VPWR VGND sg13g2_a22oi_1
X_2449_ _0739_ _0745_ _0746_ VPWR VGND sg13g2_nor2_1
XFILLER_29_525 VPWR VGND sg13g2_decap_8
X_4119_ net669 VGND VPWR net377 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[39\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_29_547 VPWR VGND sg13g2_fill_1
XFILLER_13_915 VPWR VGND sg13g2_decap_8
XFILLER_24_230 VPWR VGND sg13g2_decap_8
XFILLER_40_734 VPWR VGND sg13g2_decap_8
XFILLER_24_285 VPWR VGND sg13g2_decap_8
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_33_22 VPWR VGND sg13g2_fill_1
XFILLER_40_756 VPWR VGND sg13g2_fill_2
XFILLER_48_812 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_fill_2
XFILLER_0_885 VPWR VGND sg13g2_decap_8
Xhold7 u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[0\] VPWR VGND net49 sg13g2_dlygate4sd3_1
XFILLER_48_889 VPWR VGND sg13g2_decap_8
XFILLER_31_701 VPWR VGND sg13g2_fill_2
XFILLER_8_952 VPWR VGND sg13g2_decap_8
XFILLER_11_480 VPWR VGND sg13g2_fill_1
XFILLER_11_491 VPWR VGND sg13g2_fill_2
Xhold418 u_usb_cdc.u_sie.delay_cnt_q\[2\] VPWR VGND net460 sg13g2_dlygate4sd3_1
Xhold407 _0151_ VPWR VGND net449 sg13g2_dlygate4sd3_1
XFILLER_7_495 VPWR VGND sg13g2_fill_2
X_3421_ net778 net775 net783 _1437_ VPWR VGND _0548_ sg13g2_nand4_1
Xhold429 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[33\] VPWR VGND
+ net471 sg13g2_dlygate4sd3_1
X_3352_ VGND VPWR _1895_ net570 _0276_ _1390_ sg13g2_a21oi_1
X_2303_ _0604_ net745 net833 VPWR VGND sg13g2_nand2_2
X_3283_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[7\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[15\]
+ net818 _1348_ VPWR VGND sg13g2_mux2_1
X_2234_ net772 u_usb_cdc.u_ctrl_endp.max_length_q\[5\] _0536_ VPWR VGND sg13g2_xor2_1
X_2165_ _1922_ u_usb_cdc.u_sie.pid_q\[1\] _0467_ VPWR VGND sg13g2_nor2_1
X_2096_ VPWR _1974_ net337 VGND sg13g2_inv_1
XFILLER_22_745 VPWR VGND sg13g2_fill_1
XFILLER_10_918 VPWR VGND sg13g2_decap_8
XFILLER_16_1009 VPWR VGND sg13g2_decap_8
X_2998_ _1142_ net157 net614 VPWR VGND sg13g2_nand2_1
XFILLER_21_266 VPWR VGND sg13g2_fill_1
X_3619_ _1525_ _1549_ _0665_ _1592_ VPWR VGND sg13g2_nand3_1
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_1_638 VPWR VGND sg13g2_decap_8
XFILLER_29_311 VPWR VGND sg13g2_decap_4
XFILLER_45_804 VPWR VGND sg13g2_fill_1
XFILLER_28_33 VPWR VGND sg13g2_fill_2
XFILLER_17_506 VPWR VGND sg13g2_decap_8
XFILLER_17_517 VPWR VGND sg13g2_fill_1
XFILLER_17_528 VPWR VGND sg13g2_decap_4
XFILLER_28_77 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_fill_1
XFILLER_44_347 VPWR VGND sg13g2_fill_1
XFILLER_44_369 VPWR VGND sg13g2_decap_4
XFILLER_13_701 VPWR VGND sg13g2_decap_8
XFILLER_12_233 VPWR VGND sg13g2_decap_4
XFILLER_40_553 VPWR VGND sg13g2_decap_8
XFILLER_40_586 VPWR VGND sg13g2_fill_1
XFILLER_8_248 VPWR VGND sg13g2_fill_2
XFILLER_5_911 VPWR VGND sg13g2_decap_8
XFILLER_4_421 VPWR VGND sg13g2_fill_2
XFILLER_5_988 VPWR VGND sg13g2_decap_8
XFILLER_4_465 VPWR VGND sg13g2_fill_1
XFILLER_0_682 VPWR VGND sg13g2_decap_8
XFILLER_48_697 VPWR VGND sg13g2_fill_1
XFILLER_35_347 VPWR VGND sg13g2_fill_1
X_3970_ _1858_ u_usb_cdc.u_sie.data_q\[6\] net834 _1944_ net838 VPWR VGND sg13g2_a22oi_1
X_2921_ _1107_ VPWR _0128_ VGND _1074_ net615 sg13g2_o21ai_1
XFILLER_44_892 VPWR VGND sg13g2_decap_8
X_2852_ _1072_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2783_ u_usb_cdc.u_ctrl_endp.in_endp_q _0991_ u_usb_cdc.u_ctrl_endp.endp_q\[1\] _1027_
+ VPWR VGND sg13g2_nand3_1
Xhold204 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[41\] VPWR
+ VGND net246 sg13g2_dlygate4sd3_1
Xhold226 _0189_ VPWR VGND net268 sg13g2_dlygate4sd3_1
Xhold215 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[4\] VPWR VGND net257 sg13g2_dlygate4sd3_1
X_4453_ net672 VGND VPWR _0439_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
Xhold248 _0319_ VPWR VGND net290 sg13g2_dlygate4sd3_1
Xhold259 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[0\] VPWR VGND
+ net301 sg13g2_dlygate4sd3_1
Xhold237 _0385_ VPWR VGND net279 sg13g2_dlygate4sd3_1
X_3404_ _0647_ VPWR _1424_ VGND _0844_ _1423_ sg13g2_o21ai_1
X_4384_ net722 VGND VPWR net288 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[5\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
Xfanout706 _1986_ net706 VPWR VGND sg13g2_buf_8
X_3335_ VGND VPWR net717 net569 _0267_ _1382_ sg13g2_a21oi_1
Xfanout717 _1900_ net717 VPWR VGND sg13g2_buf_8
Xfanout739 net744 net739 VPWR VGND sg13g2_buf_8
Xfanout728 net732 net728 VPWR VGND sg13g2_buf_8
X_3266_ _0248_ _1332_ _1331_ VPWR VGND sg13g2_nand2b_1
X_2217_ _0519_ _0517_ _0518_ VPWR VGND sg13g2_nand2_1
X_3197_ _1270_ net768 net960 VPWR VGND sg13g2_nand2_1
X_2148_ _0451_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[3\] _0450_ VPWR VGND sg13g2_nand2_1
XFILLER_38_196 VPWR VGND sg13g2_fill_1
X_2079_ VPWR _1958_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[1\] VGND sg13g2_inv_1
XFILLER_34_380 VPWR VGND sg13g2_fill_1
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_1_435 VPWR VGND sg13g2_decap_8
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_9_502 VPWR VGND sg13g2_fill_1
XFILLER_13_564 VPWR VGND sg13g2_decap_4
XFILLER_13_597 VPWR VGND sg13g2_decap_8
XFILLER_5_785 VPWR VGND sg13g2_decap_8
XFILLER_4_273 VPWR VGND sg13g2_fill_2
XFILLER_45_1024 VPWR VGND sg13g2_decap_4
X_3120_ net323 net605 _1216_ VPWR VGND sg13g2_nor2_1
XFILLER_49_984 VPWR VGND sg13g2_decap_8
X_3051_ _1178_ net753 net630 VPWR VGND sg13g2_nand2_2
XFILLER_36_667 VPWR VGND sg13g2_fill_1
X_3953_ _0424_ _1841_ _1843_ net621 _1976_ VPWR VGND sg13g2_a22oi_1
XFILLER_16_380 VPWR VGND sg13g2_fill_2
XFILLER_16_391 VPWR VGND sg13g2_fill_1
X_2904_ net454 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ _1100_ _0118_ VPWR VGND sg13g2_mux2_1
X_3884_ net357 net743 _1796_ VPWR VGND sg13g2_nor2_1
X_2835_ _1039_ _1057_ net828 _1059_ VPWR VGND sg13g2_nand3_1
X_2766_ net832 _1010_ _1011_ _1012_ VPWR VGND sg13g2_nor3_1
X_2697_ net829 VPWR _0958_ VGND net622 _2003_ sg13g2_o21ai_1
X_4436_ net696 VGND VPWR _0427_ u_usb_cdc.u_sie.u_phy_tx.data_q\[6\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_4367_ net689 VGND VPWR net1019 u_usb_cdc.u_sie.pid_q\[3\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_3318_ _1358_ _1371_ _1372_ VPWR VGND sg13g2_nor2_1
Xfanout569 _1377_ net569 VPWR VGND sg13g2_buf_8
X_4298_ net674 VGND VPWR _0300_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[5\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_3249_ net816 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[36\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[44\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[52\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[60\] net811 _1317_
+ VPWR VGND sg13g2_mux4_1
XFILLER_26_188 VPWR VGND sg13g2_decap_4
XFILLER_41_55 VPWR VGND sg13g2_fill_2
XFILLER_10_556 VPWR VGND sg13g2_fill_1
XFILLER_9_2 VPWR VGND sg13g2_fill_1
XFILLER_2_711 VPWR VGND sg13g2_decap_8
Xhold590 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[7\] VPWR VGND net908 sg13g2_dlygate4sd3_1
XFILLER_49_214 VPWR VGND sg13g2_decap_4
XFILLER_2_788 VPWR VGND sg13g2_decap_8
XFILLER_1_265 VPWR VGND sg13g2_decap_4
XFILLER_46_921 VPWR VGND sg13g2_decap_8
XFILLER_18_623 VPWR VGND sg13g2_fill_1
XFILLER_46_998 VPWR VGND sg13g2_decap_8
XFILLER_14_873 VPWR VGND sg13g2_decap_4
X_2620_ _0898_ VPWR _0023_ VGND _0613_ _0894_ sg13g2_o21ai_1
X_2551_ _0722_ VPWR _0841_ VGND _0700_ _0710_ sg13g2_o21ai_1
X_2482_ VGND VPWR _0779_ _0778_ net717 sg13g2_or2_1
X_4221_ net661 VGND VPWR _0224_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[57\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_4152_ net683 VGND VPWR _0155_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[1\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_4083_ net656 VGND VPWR net408 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[3\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3103_ _1207_ net64 _1202_ VPWR VGND sg13g2_nand2_1
XFILLER_49_781 VPWR VGND sg13g2_decap_8
X_3034_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\] net709
+ _1964_ _1136_ _1166_ VPWR VGND sg13g2_and4_1
XFILLER_37_954 VPWR VGND sg13g2_decap_8
XFILLER_23_103 VPWR VGND sg13g2_fill_1
XFILLER_24_648 VPWR VGND sg13g2_fill_2
X_3936_ u_usb_cdc.ctrl_stall _0572_ net839 _1828_ VPWR VGND sg13g2_nand3_1
X_3867_ net566 _1782_ _1785_ VPWR VGND sg13g2_nor2_1
X_3798_ VPWR _0379_ _1733_ VGND sg13g2_inv_1
X_2818_ net3 net1021 net637 _0076_ VPWR VGND sg13g2_mux2_1
XFILLER_11_58 VPWR VGND sg13g2_decap_8
X_2749_ net747 _0995_ _0996_ VPWR VGND sg13g2_nor2_1
X_4419_ net730 VGND VPWR _0418_ u_usb_cdc.u_sie.rx_data\[6\] clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_28_921 VPWR VGND sg13g2_fill_2
XFILLER_28_998 VPWR VGND sg13g2_decap_8
XFILLER_43_957 VPWR VGND sg13g2_decap_8
XFILLER_42_445 VPWR VGND sg13g2_fill_2
XFILLER_42_478 VPWR VGND sg13g2_fill_1
XFILLER_30_629 VPWR VGND sg13g2_fill_2
XFILLER_11_821 VPWR VGND sg13g2_fill_2
XFILLER_11_832 VPWR VGND sg13g2_fill_2
XFILLER_23_670 VPWR VGND sg13g2_decap_8
XFILLER_7_803 VPWR VGND sg13g2_decap_8
XFILLER_22_191 VPWR VGND sg13g2_fill_2
XFILLER_10_386 VPWR VGND sg13g2_fill_2
XFILLER_42_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_585 VPWR VGND sg13g2_decap_8
XFILLER_37_239 VPWR VGND sg13g2_fill_1
XFILLER_46_795 VPWR VGND sg13g2_decap_8
XFILLER_45_272 VPWR VGND sg13g2_fill_1
XFILLER_34_924 VPWR VGND sg13g2_decap_8
XFILLER_33_478 VPWR VGND sg13g2_fill_1
X_3721_ _1686_ VPWR _0349_ VGND _1897_ net598 sg13g2_o21ai_1
X_3652_ _1622_ _1623_ _1624_ VPWR VGND sg13g2_nor2_1
X_2603_ _0467_ _0495_ net706 _0884_ VPWR VGND _0883_ sg13g2_nand4_1
X_3583_ VGND VPWR _1541_ _1556_ _1558_ _1557_ sg13g2_a21oi_1
XFILLER_6_891 VPWR VGND sg13g2_decap_8
X_2534_ _0828_ net717 _0698_ VPWR VGND sg13g2_nand2_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_2465_ _0714_ _0747_ _0675_ _0762_ VPWR VGND sg13g2_nand3_1
X_4204_ net659 VGND VPWR net79 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[40\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_2396_ net586 net584 net619 _0686_ _0696_ VPWR VGND sg13g2_nor4_1
XFILLER_3_92 VPWR VGND sg13g2_fill_1
X_4135_ net670 VGND VPWR net60 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[55\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_28_206 VPWR VGND sg13g2_decap_4
X_4066_ net698 VGND VPWR net558 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
X_3017_ net823 _1150_ net756 _1155_ VPWR VGND sg13g2_nand3_1
XFILLER_24_401 VPWR VGND sg13g2_decap_4
XFILLER_24_478 VPWR VGND sg13g2_fill_2
XFILLER_40_949 VPWR VGND sg13g2_decap_8
X_3919_ _1812_ VPWR _1813_ VGND net282 net705 sg13g2_o21ai_1
XFILLER_47_515 VPWR VGND sg13g2_decap_8
XFILLER_27_283 VPWR VGND sg13g2_fill_1
XFILLER_42_253 VPWR VGND sg13g2_fill_1
XFILLER_31_916 VPWR VGND sg13g2_fill_1
XFILLER_11_651 VPWR VGND sg13g2_fill_2
XFILLER_10_161 VPWR VGND sg13g2_fill_2
XFILLER_7_611 VPWR VGND sg13g2_fill_2
XFILLER_3_850 VPWR VGND sg13g2_decap_8
XFILLER_2_371 VPWR VGND sg13g2_decap_8
X_2250_ net773 net770 _0552_ VPWR VGND sg13g2_nor2_2
X_2181_ _0483_ _0481_ _0482_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_773 VPWR VGND sg13g2_fill_1
X_3704_ net794 VPWR _1673_ VGND net801 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[55\]
+ sg13g2_o21ai_1
X_3635_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[20\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[28\]
+ net801 _1607_ VPWR VGND sg13g2_mux2_1
X_3566_ VGND VPWR net631 _1540_ _1541_ _1489_ sg13g2_a21oi_1
X_3497_ _0326_ net572 _0503_ net575 _1948_ VPWR VGND sg13g2_a22oi_1
X_2517_ _0813_ _0698_ _0713_ VPWR VGND sg13g2_nand2_1
X_2448_ u_usb_cdc.sie_out_data\[5\] net717 u_usb_cdc.configured_o _0744_ _0745_ VPWR
+ VGND sg13g2_and4_1
X_2379_ net586 net583 _0653_ net619 _0679_ VPWR VGND sg13g2_nor4_1
X_4118_ net670 VGND VPWR net476 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[38\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_44_529 VPWR VGND sg13g2_fill_2
X_4049_ net694 VGND VPWR net187 u_usb_cdc.u_sie.phy_state_q\[5\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_40_713 VPWR VGND sg13g2_decap_8
XFILLER_25_787 VPWR VGND sg13g2_fill_1
XFILLER_4_669 VPWR VGND sg13g2_decap_8
XFILLER_0_864 VPWR VGND sg13g2_decap_8
Xhold8 _0046_ VPWR VGND net50 sg13g2_dlygate4sd3_1
XFILLER_48_868 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_35_518 VPWR VGND sg13g2_fill_2
XFILLER_31_713 VPWR VGND sg13g2_fill_1
XFILLER_8_931 VPWR VGND sg13g2_decap_8
XFILLER_7_441 VPWR VGND sg13g2_fill_1
XFILLER_12_993 VPWR VGND sg13g2_decap_8
Xhold408 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[64\] VPWR VGND
+ net450 sg13g2_dlygate4sd3_1
Xhold419 _0318_ VPWR VGND net461 sg13g2_dlygate4sd3_1
X_3420_ _1436_ net775 _1424_ VPWR VGND sg13g2_nand2_1
XFILLER_48_1022 VPWR VGND sg13g2_decap_8
X_3351_ net391 net570 _1390_ VPWR VGND sg13g2_nor2_1
X_2302_ _0603_ net745 _1904_ VPWR VGND sg13g2_nand2_1
X_3282_ _1278_ _1345_ _1346_ _1347_ VPWR VGND sg13g2_nor3_1
XFILLER_39_802 VPWR VGND sg13g2_fill_1
X_2233_ u_usb_cdc.u_ctrl_endp.max_length_q\[4\] net775 _0535_ VPWR VGND sg13g2_xor2_1
XFILLER_39_824 VPWR VGND sg13g2_decap_4
X_2164_ _0459_ _0463_ _0458_ _0466_ VPWR VGND _0465_ sg13g2_nand4_1
X_2095_ VPWR _1973_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[15\]
+ VGND sg13g2_inv_1
XFILLER_34_584 VPWR VGND sg13g2_fill_2
X_2997_ _1141_ VPWR _0170_ VGND net719 net614 sg13g2_o21ai_1
X_3618_ _1583_ VPWR _1591_ VGND net788 _1590_ sg13g2_o21ai_1
XFILLER_1_617 VPWR VGND sg13g2_decap_8
X_3549_ net774 _1918_ _1525_ VPWR VGND sg13g2_nor2_1
XFILLER_45_849 VPWR VGND sg13g2_decap_8
XFILLER_5_967 VPWR VGND sg13g2_decap_8
XFILLER_0_661 VPWR VGND sg13g2_decap_8
XFILLER_44_871 VPWR VGND sg13g2_decap_8
X_2920_ _1107_ net56 _1101_ VPWR VGND sg13g2_nand2_1
XFILLER_43_392 VPWR VGND sg13g2_fill_1
XFILLER_31_521 VPWR VGND sg13g2_decap_8
XFILLER_31_532 VPWR VGND sg13g2_fill_1
XFILLER_31_587 VPWR VGND sg13g2_decap_8
X_2851_ _1071_ net69 _1059_ VPWR VGND sg13g2_nand2_1
X_2782_ _1987_ _1020_ u_usb_cdc.endp\[1\] _1026_ VPWR VGND sg13g2_nand3_1
XFILLER_8_783 VPWR VGND sg13g2_decap_8
X_4452_ net683 VGND VPWR _0438_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
Xhold205 _0208_ VPWR VGND net247 sg13g2_dlygate4sd3_1
Xhold216 _0032_ VPWR VGND net258 sg13g2_dlygate4sd3_1
Xhold238 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[2\] VPWR VGND
+ net280 sg13g2_dlygate4sd3_1
Xhold227 u_usb_cdc.u_ctrl_endp.addr_dd\[0\] VPWR VGND net269 sg13g2_dlygate4sd3_1
Xhold249 u_usb_cdc.u_sie.out_eop_q VPWR VGND net291 sg13g2_dlygate4sd3_1
X_3403_ u_usb_cdc.u_ctrl_endp.state_q\[3\] _1422_ _1423_ VPWR VGND sg13g2_nor2_1
X_4383_ net722 VGND VPWR net279 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[4\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
Xfanout707 _1965_ net707 VPWR VGND sg13g2_buf_8
X_3334_ net479 _1377_ _1382_ VPWR VGND sg13g2_nor2_1
Xfanout718 _1897_ net718 VPWR VGND sg13g2_buf_8
Xfanout729 net732 net729 VPWR VGND sg13g2_buf_8
X_3265_ _1332_ _1296_ net134 net602 net897 VPWR VGND sg13g2_a22oi_1
X_2216_ _0518_ _0504_ _0509_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_1025 VPWR VGND sg13g2_decap_4
X_3196_ _1269_ _0735_ _1250_ VPWR VGND sg13g2_nand2_1
XFILLER_27_827 VPWR VGND sg13g2_fill_2
XFILLER_38_164 VPWR VGND sg13g2_fill_2
X_2147_ _1937_ net703 _0450_ VPWR VGND sg13g2_nor2_2
XFILLER_26_337 VPWR VGND sg13g2_fill_1
X_2078_ VPWR _1957_ net525 VGND sg13g2_inv_1
XFILLER_10_738 VPWR VGND sg13g2_fill_2
XFILLER_6_709 VPWR VGND sg13g2_decap_8
XFILLER_30_35 VPWR VGND sg13g2_decap_8
XFILLER_1_414 VPWR VGND sg13g2_decap_8
Xhold750 u_usb_cdc.sie_out_err VPWR VGND net1068 sg13g2_dlygate4sd3_1
XFILLER_44_178 VPWR VGND sg13g2_fill_1
XFILLER_41_841 VPWR VGND sg13g2_fill_1
XFILLER_40_362 VPWR VGND sg13g2_decap_8
XFILLER_13_587 VPWR VGND sg13g2_decap_8
XFILLER_5_764 VPWR VGND sg13g2_decap_8
XFILLER_45_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_296 VPWR VGND sg13g2_fill_1
XFILLER_1_981 VPWR VGND sg13g2_decap_8
X_3050_ net283 net612 _1177_ VPWR VGND sg13g2_nor2_1
XFILLER_49_963 VPWR VGND sg13g2_decap_8
XFILLER_48_495 VPWR VGND sg13g2_decap_8
XFILLER_35_112 VPWR VGND sg13g2_decap_4
XFILLER_17_871 VPWR VGND sg13g2_decap_8
X_3952_ VGND VPWR u_usb_cdc.u_sie.u_phy_tx.data_q\[4\] _1842_ _1843_ net621 sg13g2_a21oi_1
XFILLER_32_852 VPWR VGND sg13g2_decap_4
X_2903_ net446 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ _1100_ _0117_ VPWR VGND sg13g2_mux2_1
X_3883_ _1794_ _1795_ _0402_ VPWR VGND sg13g2_nor2_1
X_2834_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ net438 _1058_ _0090_ VPWR VGND sg13g2_mux2_1
XFILLER_31_373 VPWR VGND sg13g2_fill_2
XFILLER_32_896 VPWR VGND sg13g2_fill_1
X_2765_ _1011_ _1966_ net634 VPWR VGND sg13g2_xnor2_1
X_2696_ _0957_ net556 _0953_ VPWR VGND sg13g2_nand2_1
X_4435_ net696 VGND VPWR net275 u_usb_cdc.u_sie.u_phy_tx.data_q\[5\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_6_81 VPWR VGND sg13g2_fill_1
X_4366_ net694 VGND VPWR net1010 u_usb_cdc.u_sie.pid_q\[2\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3317_ net280 _1370_ _1128_ _1371_ VPWR VGND sg13g2_mux2_1
X_4297_ net674 VGND VPWR _0299_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[4\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
X_3248_ _0246_ _1316_ _1315_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_462 VPWR VGND sg13g2_fill_1
X_3179_ _1255_ _0735_ _1240_ VPWR VGND sg13g2_nand2_1
XFILLER_26_101 VPWR VGND sg13g2_decap_4
XFILLER_26_134 VPWR VGND sg13g2_decap_4
XFILLER_26_167 VPWR VGND sg13g2_decap_4
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_25_79 VPWR VGND sg13g2_fill_2
XFILLER_23_885 VPWR VGND sg13g2_fill_1
XFILLER_2_767 VPWR VGND sg13g2_decap_8
Xhold580 _0248_ VPWR VGND net898 sg13g2_dlygate4sd3_1
Xhold591 _1727_ VPWR VGND net909 sg13g2_dlygate4sd3_1
XFILLER_46_900 VPWR VGND sg13g2_decap_8
XFILLER_46_977 VPWR VGND sg13g2_decap_8
XFILLER_18_646 VPWR VGND sg13g2_decap_8
XFILLER_32_126 VPWR VGND sg13g2_decap_8
XFILLER_41_660 VPWR VGND sg13g2_decap_8
XFILLER_41_682 VPWR VGND sg13g2_decap_4
XFILLER_14_896 VPWR VGND sg13g2_fill_1
XFILLER_9_355 VPWR VGND sg13g2_fill_1
X_2550_ _0719_ _0823_ _0718_ _0840_ VPWR VGND sg13g2_nand3_1
X_2481_ u_usb_cdc.u_ctrl_endp.req_q\[7\] _0688_ net738 _0778_ VPWR VGND sg13g2_nand3_1
XFILLER_49_4 VPWR VGND sg13g2_decap_8
X_4220_ net665 VGND VPWR net224 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[56\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_4151_ net674 VGND VPWR net492 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[71\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_49_760 VPWR VGND sg13g2_decap_8
X_4082_ net651 VGND VPWR net425 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[2\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3102_ _1206_ VPWR _0210_ VGND net708 _1157_ sg13g2_o21ai_1
X_3033_ _1164_ VPWR _0182_ VGND u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[2\]
+ _1165_ sg13g2_o21ai_1
XFILLER_37_933 VPWR VGND sg13g2_decap_8
XFILLER_36_454 VPWR VGND sg13g2_fill_2
XFILLER_24_627 VPWR VGND sg13g2_decap_8
X_3935_ _1827_ net211 net621 VPWR VGND sg13g2_nand2_1
XFILLER_32_693 VPWR VGND sg13g2_decap_4
X_3866_ _1784_ net711 net566 VPWR VGND sg13g2_nand2_1
X_3797_ _1733_ _1719_ _1732_ net579 net908 VPWR VGND sg13g2_a22oi_1
X_2817_ net2 net1022 net637 _0075_ VPWR VGND sg13g2_mux2_1
X_2748_ _0994_ _0990_ _0995_ VPWR VGND sg13g2_nor2b_1
X_2679_ _0440_ net635 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] _0946_ VPWR VGND sg13g2_nand3_1
X_4418_ net730 VGND VPWR _0417_ u_usb_cdc.u_sie.rx_data\[5\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_4349_ net681 VGND VPWR _0351_ u_usb_cdc.sie_out_data\[4\] clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_28_977 VPWR VGND sg13g2_decap_8
XFILLER_43_936 VPWR VGND sg13g2_decap_8
XFILLER_27_465 VPWR VGND sg13g2_decap_4
XFILLER_35_1013 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_fill_2
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_38_719 VPWR VGND sg13g2_fill_1
XFILLER_37_207 VPWR VGND sg13g2_fill_2
XFILLER_46_774 VPWR VGND sg13g2_decap_8
XFILLER_42_991 VPWR VGND sg13g2_decap_8
X_3720_ net591 _1683_ net762 _1686_ VPWR VGND sg13g2_nand3_1
XFILLER_13_181 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_40_clk clknet_3_5__leaf_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_3651_ net625 VPWR _1623_ VGND _0576_ _1615_ sg13g2_o21ai_1
X_2602_ VGND VPWR _1924_ u_usb_cdc.u_sie.pid_q\[3\] _0883_ net762 sg13g2_a21oi_1
X_3582_ net597 VPWR _1557_ VGND net940 net624 sg13g2_o21ai_1
XFILLER_6_870 VPWR VGND sg13g2_decap_8
X_2533_ _0826_ VPWR _0007_ VGND _0741_ _0827_ sg13g2_o21ai_1
X_2464_ VGND VPWR _0759_ _0760_ _0761_ net617 sg13g2_a21oi_1
X_4203_ net662 VGND VPWR net142 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[39\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2395_ net587 net584 net620 _0695_ VPWR VGND sg13g2_nor3_2
X_4134_ net670 VGND VPWR net88 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[54\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_3_1011 VPWR VGND sg13g2_decap_8
X_4065_ net698 VGND VPWR net932 _0053_ clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3016_ _1154_ net122 _1146_ VPWR VGND sg13g2_nand2_1
XFILLER_36_262 VPWR VGND sg13g2_fill_2
XFILLER_25_958 VPWR VGND sg13g2_decap_8
XFILLER_25_969 VPWR VGND sg13g2_fill_1
XFILLER_36_295 VPWR VGND sg13g2_fill_1
XFILLER_40_928 VPWR VGND sg13g2_decap_8
XFILLER_11_118 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_31_clk clknet_3_7__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_3918_ _1811_ _1808_ _1807_ _1812_ VPWR VGND sg13g2_a21o_1
X_3849_ _1770_ VPWR _0392_ VGND _1740_ _1771_ sg13g2_o21ai_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_229 VPWR VGND sg13g2_fill_2
XFILLER_28_774 VPWR VGND sg13g2_fill_2
XFILLER_16_969 VPWR VGND sg13g2_fill_1
XFILLER_31_906 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_22_clk clknet_3_3__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_7_689 VPWR VGND sg13g2_fill_1
XFILLER_12_91 VPWR VGND sg13g2_fill_2
XFILLER_40_8 VPWR VGND sg13g2_fill_2
X_2180_ _0482_ u_usb_cdc.sie_out_data\[3\] net752 VPWR VGND sg13g2_xnor2_1
XFILLER_18_251 VPWR VGND sg13g2_fill_1
XFILLER_46_571 VPWR VGND sg13g2_fill_1
XFILLER_34_766 VPWR VGND sg13g2_decap_8
XFILLER_21_427 VPWR VGND sg13g2_decap_4
XFILLER_33_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_3703_ VGND VPWR net802 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[47\]
+ _1672_ _1671_ sg13g2_a21oi_1
X_3634_ VGND VPWR net799 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[12\]
+ _1606_ _1605_ sg13g2_a21oi_1
X_3565_ _1532_ VPWR _1540_ VGND net788 _1539_ sg13g2_o21ai_1
X_3496_ _0325_ net572 _0520_ net575 _1949_ VPWR VGND sg13g2_a22oi_1
X_2516_ _0809_ _0812_ _0742_ _0004_ VPWR VGND sg13g2_nand3_1
X_2447_ net755 net756 u_usb_cdc.sie_out_data\[4\] net752 _0744_ VPWR VGND sg13g2_nor4_1
XFILLER_25_1012 VPWR VGND sg13g2_decap_8
X_2378_ VGND VPWR _0659_ _0674_ _0678_ _0677_ sg13g2_a21oi_1
X_4117_ net655 VGND VPWR net514 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[37\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_4048_ net687 VGND VPWR _0023_ u_usb_cdc.u_sie.phy_state_q\[4\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_37_571 VPWR VGND sg13g2_decap_8
XFILLER_24_265 VPWR VGND sg13g2_decap_8
XFILLER_12_449 VPWR VGND sg13g2_decap_8
XFILLER_32_1027 VPWR VGND sg13g2_fill_2
XFILLER_4_604 VPWR VGND sg13g2_decap_8
XFILLER_4_648 VPWR VGND sg13g2_decap_8
XFILLER_3_103 VPWR VGND sg13g2_fill_2
XFILLER_0_843 VPWR VGND sg13g2_decap_8
Xhold9 u_usb_cdc.clk_cnt_q\[1\] VPWR VGND net51 sg13g2_dlygate4sd3_1
XFILLER_48_847 VPWR VGND sg13g2_decap_8
XFILLER_47_324 VPWR VGND sg13g2_fill_1
XFILLER_16_700 VPWR VGND sg13g2_decap_8
XFILLER_31_703 VPWR VGND sg13g2_fill_1
XFILLER_43_563 VPWR VGND sg13g2_decap_8
XFILLER_8_910 VPWR VGND sg13g2_decap_8
XFILLER_12_972 VPWR VGND sg13g2_decap_8
XFILLER_11_493 VPWR VGND sg13g2_fill_1
XFILLER_8_987 VPWR VGND sg13g2_decap_8
Xhold409 _0147_ VPWR VGND net451 sg13g2_dlygate4sd3_1
XFILLER_48_1001 VPWR VGND sg13g2_decap_8
X_3350_ VGND VPWR _1894_ net570 _0275_ _1389_ sg13g2_a21oi_1
X_2301_ _0597_ VPWR _0063_ VGND _0531_ net261 sg13g2_o21ai_1
X_3281_ net201 net818 _1346_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_4 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_2_clk clknet_3_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_2232_ net785 u_usb_cdc.u_ctrl_endp.max_length_q\[1\] _0534_ VPWR VGND sg13g2_xor2_1
X_2163_ _0460_ _0461_ _0462_ _0464_ _0465_ VPWR VGND sg13g2_nor4_1
XFILLER_47_891 VPWR VGND sg13g2_decap_8
X_2094_ VPWR _1972_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[45\]
+ VGND sg13g2_inv_1
XFILLER_0_1025 VPWR VGND sg13g2_decap_4
XFILLER_34_530 VPWR VGND sg13g2_fill_1
XFILLER_34_596 VPWR VGND sg13g2_decap_8
X_2996_ _1141_ net63 net614 VPWR VGND sg13g2_nand2_1
X_3617_ _1589_ VPWR _1590_ VGND net789 _1584_ sg13g2_o21ai_1
X_3548_ _1504_ _1507_ net776 _1524_ VPWR VGND sg13g2_nand3_1
X_3479_ _1474_ net319 net594 VPWR VGND sg13g2_nand2_1
XFILLER_45_828 VPWR VGND sg13g2_decap_8
XFILLER_29_357 VPWR VGND sg13g2_decap_8
XFILLER_29_368 VPWR VGND sg13g2_fill_2
XFILLER_44_67 VPWR VGND sg13g2_fill_2
XFILLER_9_718 VPWR VGND sg13g2_fill_2
XFILLER_8_228 VPWR VGND sg13g2_decap_8
XFILLER_5_946 VPWR VGND sg13g2_decap_8
XFILLER_0_640 VPWR VGND sg13g2_decap_8
XFILLER_48_666 VPWR VGND sg13g2_fill_2
XFILLER_48_655 VPWR VGND sg13g2_decap_8
XFILLER_44_850 VPWR VGND sg13g2_decap_8
XFILLER_16_552 VPWR VGND sg13g2_fill_1
XFILLER_18_90 VPWR VGND sg13g2_fill_1
XFILLER_31_500 VPWR VGND sg13g2_decap_8
X_2850_ _1069_ VPWR _0094_ VGND net616 _1070_ sg13g2_o21ai_1
XFILLER_43_382 VPWR VGND sg13g2_fill_1
X_2781_ _1025_ net354 _1024_ VPWR VGND sg13g2_nand2_1
XFILLER_8_762 VPWR VGND sg13g2_decap_8
Xhold206 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[60\] VPWR
+ VGND net248 sg13g2_dlygate4sd3_1
Xhold217 u_usb_cdc.u_sie.phy_state_q\[10\] VPWR VGND net259 sg13g2_dlygate4sd3_1
X_4451_ net684 VGND VPWR net166 u_usb_cdc.u_sie.in_zlp_q\[0\] clknet_leaf_25_clk sg13g2_dfrbpq_1
Xhold239 _0165_ VPWR VGND net281 sg13g2_dlygate4sd3_1
Xhold228 _0268_ VPWR VGND net270 sg13g2_dlygate4sd3_1
XFILLER_7_294 VPWR VGND sg13g2_decap_4
X_3402_ VGND VPWR _0554_ _0640_ _1422_ _1920_ sg13g2_a21oi_1
X_4382_ net722 VGND VPWR net1008 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[3\] clknet_leaf_46_clk
+ sg13g2_dfrbpq_1
X_3333_ VGND VPWR net719 net569 _0266_ _1381_ sg13g2_a21oi_1
Xfanout719 _1896_ net719 VPWR VGND sg13g2_buf_8
Xfanout708 _1963_ net708 VPWR VGND sg13g2_buf_8
X_3264_ net805 net602 _1330_ _1331_ VPWR VGND sg13g2_nor3_1
XFILLER_22_0 VPWR VGND sg13g2_fill_1
X_2215_ _0517_ net918 _0510_ VPWR VGND sg13g2_xnor2_1
X_3195_ _1254_ net820 _1268_ _0241_ VPWR VGND sg13g2_a21o_1
X_2146_ _0449_ net49 net521 VPWR VGND sg13g2_nand2b_1
X_2077_ VPWR _1956_ net186 VGND sg13g2_inv_1
XFILLER_10_706 VPWR VGND sg13g2_decap_4
X_2979_ _1131_ net301 _1130_ VPWR VGND sg13g2_nand2_1
XFILLER_2_949 VPWR VGND sg13g2_decap_8
Xhold751 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\] VPWR
+ VGND net1069 sg13g2_dlygate4sd3_1
Xhold740 _0241_ VPWR VGND net1058 sg13g2_dlygate4sd3_1
XFILLER_39_12 VPWR VGND sg13g2_decap_4
XFILLER_17_338 VPWR VGND sg13g2_fill_1
XFILLER_25_360 VPWR VGND sg13g2_fill_1
XFILLER_13_544 VPWR VGND sg13g2_decap_8
XFILLER_25_393 VPWR VGND sg13g2_fill_2
XFILLER_40_341 VPWR VGND sg13g2_decap_8
XFILLER_9_548 VPWR VGND sg13g2_fill_2
XFILLER_5_743 VPWR VGND sg13g2_decap_8
XFILLER_1_960 VPWR VGND sg13g2_decap_8
XFILLER_49_942 VPWR VGND sg13g2_decap_8
XFILLER_35_135 VPWR VGND sg13g2_fill_2
X_3951_ _1805_ VPWR _1842_ VGND _1994_ _1034_ sg13g2_o21ai_1
XFILLER_23_319 VPWR VGND sg13g2_fill_2
X_2902_ net471 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ _1100_ _0116_ VPWR VGND sg13g2_mux2_1
X_3882_ VGND VPWR net742 net287 _1795_ net878 sg13g2_a21oi_1
XFILLER_31_352 VPWR VGND sg13g2_fill_2
X_2833_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net380 _1058_ _0089_ VPWR VGND sg13g2_mux2_1
X_2764_ _0980_ _1009_ net591 _1010_ VPWR VGND sg13g2_nand3_1
X_2695_ _0956_ VPWR _0037_ VGND net382 _2000_ sg13g2_o21ai_1
X_4434_ net698 VGND VPWR _0425_ u_usb_cdc.u_sie.u_phy_tx.data_q\[4\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_4365_ net695 VGND VPWR _0367_ u_usb_cdc.u_sie.pid_q\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3316_ _1368_ _1369_ _1370_ VPWR VGND sg13g2_and2_1
X_4296_ net674 VGND VPWR _0298_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[3\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_3247_ _1316_ _1296_ net193 net601 net559 VPWR VGND sg13g2_a22oi_1
X_3178_ _1254_ _1253_ _1239_ VPWR VGND sg13g2_nand2b_1
X_2129_ _2006_ VPWR _2007_ VGND _1911_ _2003_ sg13g2_o21ai_1
XFILLER_22_341 VPWR VGND sg13g2_fill_1
XFILLER_10_525 VPWR VGND sg13g2_fill_2
XFILLER_10_547 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_fill_1
XFILLER_1_201 VPWR VGND sg13g2_fill_1
XFILLER_2_746 VPWR VGND sg13g2_decap_8
Xhold581 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\] VPWR VGND net899 sg13g2_dlygate4sd3_1
Xhold570 u_usb_cdc.u_ctrl_endp.state_q\[7\] VPWR VGND net888 sg13g2_dlygate4sd3_1
Xhold592 u_usb_cdc.u_ctrl_endp.rec_q\[1\] VPWR VGND net910 sg13g2_dlygate4sd3_1
XFILLER_49_238 VPWR VGND sg13g2_fill_2
XFILLER_46_956 VPWR VGND sg13g2_decap_8
XFILLER_45_422 VPWR VGND sg13g2_decap_4
XFILLER_18_658 VPWR VGND sg13g2_decap_8
XFILLER_18_669 VPWR VGND sg13g2_fill_1
XFILLER_14_831 VPWR VGND sg13g2_fill_1
XFILLER_13_363 VPWR VGND sg13g2_decap_8
XFILLER_12_1014 VPWR VGND sg13g2_decap_8
X_2480_ _0777_ _0776_ _0739_ VPWR VGND sg13g2_nand2b_1
X_4150_ net674 VGND VPWR net470 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[70\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3101_ _1206_ net195 _1202_ VPWR VGND sg13g2_nand2_1
X_4081_ net649 VGND VPWR net443 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[1\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_3032_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[0\] _1150_
+ net751 _1165_ VPWR VGND sg13g2_nand3_1
XFILLER_37_989 VPWR VGND sg13g2_decap_8
XFILLER_23_116 VPWR VGND sg13g2_fill_2
X_3934_ _1816_ VPWR _0422_ VGND _1823_ _1826_ sg13g2_o21ai_1
X_3865_ _1781_ VPWR _0396_ VGND _1782_ _1783_ sg13g2_o21ai_1
X_2816_ _0074_ net638 _1056_ VPWR VGND sg13g2_nand2_1
X_3796_ _1731_ VPWR _1732_ VGND net360 _0942_ sg13g2_o21ai_1
X_2747_ VGND VPWR _1955_ _0993_ _0994_ net842 sg13g2_a21oi_1
X_2678_ _0945_ net257 net703 VPWR VGND sg13g2_nand2_1
X_4417_ net730 VGND VPWR net930 u_usb_cdc.u_sie.rx_data\[4\] clknet_leaf_31_clk sg13g2_dfrbpq_2
X_4348_ net681 VGND VPWR _0350_ u_usb_cdc.sie_out_data\[3\] clknet_leaf_47_clk sg13g2_dfrbpq_2
XFILLER_47_709 VPWR VGND sg13g2_decap_8
X_4279_ net680 VGND VPWR net365 u_usb_cdc.u_ctrl_endp.addr_dd\[6\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
XFILLER_27_422 VPWR VGND sg13g2_decap_8
XFILLER_28_956 VPWR VGND sg13g2_decap_8
XFILLER_43_915 VPWR VGND sg13g2_decap_8
XFILLER_15_617 VPWR VGND sg13g2_decap_8
XFILLER_14_127 VPWR VGND sg13g2_decap_4
XFILLER_42_447 VPWR VGND sg13g2_fill_1
XFILLER_23_650 VPWR VGND sg13g2_fill_2
XFILLER_22_193 VPWR VGND sg13g2_fill_1
XFILLER_2_543 VPWR VGND sg13g2_decap_8
XFILLER_46_753 VPWR VGND sg13g2_decap_8
XFILLER_18_444 VPWR VGND sg13g2_decap_4
XFILLER_34_959 VPWR VGND sg13g2_decap_8
XFILLER_26_90 VPWR VGND sg13g2_fill_1
XFILLER_42_970 VPWR VGND sg13g2_decap_8
X_3650_ _1529_ _1621_ _1622_ VPWR VGND sg13g2_nor2_1
X_2601_ _0877_ _0879_ _0875_ _0882_ VPWR VGND _0881_ sg13g2_nand4_1
X_3581_ _1528_ VPWR _1556_ VGND _1553_ _1555_ sg13g2_o21ai_1
X_2532_ _0827_ _0713_ _0803_ VPWR VGND sg13g2_nand2_1
XFILLER_5_381 VPWR VGND sg13g2_decap_8
X_4202_ net644 VGND VPWR net140 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[38\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2463_ VGND VPWR _0662_ _0754_ _0760_ _0757_ sg13g2_a21oi_1
X_2394_ net586 net583 net620 _0673_ _0694_ VPWR VGND sg13g2_nor4_1
X_4133_ net651 VGND VPWR net107 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[53\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_29_709 VPWR VGND sg13g2_fill_2
X_4064_ net724 VGND VPWR _0035_ u_usb_cdc.u_sie.u_phy_rx.state_q\[3\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_49_591 VPWR VGND sg13g2_decap_8
X_3015_ _1152_ VPWR _0176_ VGND net821 _1153_ sg13g2_o21ai_1
XFILLER_37_731 VPWR VGND sg13g2_decap_8
XFILLER_37_775 VPWR VGND sg13g2_fill_2
XFILLER_19_1009 VPWR VGND sg13g2_decap_8
XFILLER_24_425 VPWR VGND sg13g2_fill_2
XFILLER_40_907 VPWR VGND sg13g2_decap_8
XFILLER_12_609 VPWR VGND sg13g2_decap_4
X_3917_ _1809_ _1810_ _1696_ _1811_ VPWR VGND sg13g2_nand3_1
X_3848_ _1771_ net422 _1768_ VPWR VGND sg13g2_xnor2_1
X_3779_ VPWR _0372_ net532 VGND sg13g2_inv_1
XFILLER_15_414 VPWR VGND sg13g2_fill_2
XFILLER_42_244 VPWR VGND sg13g2_decap_8
XFILLER_15_458 VPWR VGND sg13g2_fill_2
XFILLER_30_417 VPWR VGND sg13g2_decap_8
XFILLER_42_299 VPWR VGND sg13g2_decap_4
XFILLER_8_28 VPWR VGND sg13g2_fill_2
XFILLER_23_491 VPWR VGND sg13g2_fill_2
XFILLER_7_613 VPWR VGND sg13g2_fill_1
XFILLER_11_653 VPWR VGND sg13g2_fill_1
XFILLER_3_885 VPWR VGND sg13g2_decap_8
XFILLER_34_712 VPWR VGND sg13g2_decap_4
XFILLER_21_417 VPWR VGND sg13g2_decap_4
XFILLER_34_789 VPWR VGND sg13g2_fill_2
X_3702_ net801 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[39\] _1671_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_30_984 VPWR VGND sg13g2_decap_8
X_3633_ net800 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[4\] _1605_
+ VPWR VGND sg13g2_nor2b_1
X_3564_ _1538_ VPWR _1539_ VGND net789 _1533_ sg13g2_o21ai_1
X_3495_ _0324_ net573 _0514_ net576 _1947_ VPWR VGND sg13g2_a22oi_1
X_2515_ VGND VPWR _0746_ _0811_ _0812_ _0810_ sg13g2_a21oi_1
X_2446_ _0480_ _0708_ _0743_ VPWR VGND sg13g2_nor2_2
X_2377_ net586 net584 net620 _0676_ _0677_ VPWR VGND sg13g2_nor4_1
X_4116_ net668 VGND VPWR net468 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[36\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
X_4047_ net694 VGND VPWR net526 u_usb_cdc.u_sie.phy_state_q\[3\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
XFILLER_37_550 VPWR VGND sg13g2_fill_2
XFILLER_25_734 VPWR VGND sg13g2_decap_8
XFILLER_12_417 VPWR VGND sg13g2_fill_1
XFILLER_13_929 VPWR VGND sg13g2_decap_8
XFILLER_24_299 VPWR VGND sg13g2_decap_4
XFILLER_32_1006 VPWR VGND sg13g2_decap_8
XFILLER_20_472 VPWR VGND sg13g2_fill_1
XFILLER_0_822 VPWR VGND sg13g2_decap_8
XFILLER_48_826 VPWR VGND sg13g2_decap_8
XFILLER_0_899 VPWR VGND sg13g2_decap_8
XFILLER_28_550 VPWR VGND sg13g2_decap_4
XFILLER_15_222 VPWR VGND sg13g2_decap_4
XFILLER_15_266 VPWR VGND sg13g2_fill_2
XFILLER_11_450 VPWR VGND sg13g2_decap_8
XFILLER_12_951 VPWR VGND sg13g2_decap_8
XFILLER_8_966 VPWR VGND sg13g2_decap_8
XFILLER_11_461 VPWR VGND sg13g2_fill_1
XFILLER_3_682 VPWR VGND sg13g2_decap_8
X_3280_ net819 net314 _1345_ VPWR VGND sg13g2_nor2_1
X_2300_ _0497_ net591 _0494_ _0602_ VPWR VGND _0601_ sg13g2_nand4_1
X_2231_ net779 u_usb_cdc.u_ctrl_endp.max_length_q\[3\] _0533_ VPWR VGND sg13g2_xor2_1
X_2162_ u_usb_cdc.addr\[2\] net756 _0464_ VPWR VGND sg13g2_xor2_1
X_2093_ VPWR _1971_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[44\]
+ VGND sg13g2_inv_1
XFILLER_47_870 VPWR VGND sg13g2_decap_8
XFILLER_0_1004 VPWR VGND sg13g2_decap_8
XFILLER_19_583 VPWR VGND sg13g2_decap_8
XFILLER_46_380 VPWR VGND sg13g2_decap_8
XFILLER_21_203 VPWR VGND sg13g2_fill_2
XFILLER_34_586 VPWR VGND sg13g2_fill_1
X_2995_ _1140_ VPWR _0169_ VGND net718 net614 sg13g2_o21ai_1
X_3616_ _1589_ _1586_ _1588_ VPWR VGND sg13g2_nand2_1
X_3547_ _1523_ _1519_ u_usb_cdc.u_ctrl_endp.req_q\[2\] u_usb_cdc.configured_o u_usb_cdc.u_ctrl_endp.req_q\[4\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_0_107 VPWR VGND sg13g2_decap_4
X_3478_ _1473_ VPWR _0319_ VGND net289 _0894_ sg13g2_o21ai_1
X_2429_ _0727_ u_usb_cdc.u_ctrl_endp.in_dir_q _0726_ VPWR VGND sg13g2_nand2_1
XFILLER_29_347 VPWR VGND sg13g2_fill_1
XFILLER_25_520 VPWR VGND sg13g2_fill_2
XFILLER_13_715 VPWR VGND sg13g2_decap_8
XFILLER_25_564 VPWR VGND sg13g2_decap_8
XFILLER_44_79 VPWR VGND sg13g2_fill_1
XFILLER_13_748 VPWR VGND sg13g2_fill_2
XFILLER_12_247 VPWR VGND sg13g2_decap_8
XFILLER_5_925 VPWR VGND sg13g2_decap_8
XFILLER_0_696 VPWR VGND sg13g2_decap_8
XFILLER_18_80 VPWR VGND sg13g2_fill_1
XFILLER_31_545 VPWR VGND sg13g2_decap_8
XFILLER_15_1012 VPWR VGND sg13g2_decap_8
X_2780_ _1024_ _1014_ _1016_ VPWR VGND sg13g2_nand2_1
Xhold207 _0227_ VPWR VGND net249 sg13g2_dlygate4sd3_1
X_4450_ net684 VGND VPWR net86 u_usb_cdc.u_sie.in_zlp_q\[1\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_4381_ net722 VGND VPWR net203 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[2\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_2
Xhold229 u_usb_cdc.u_ctrl_endp.endp_q\[3\] VPWR VGND net271 sg13g2_dlygate4sd3_1
X_3401_ VGND VPWR net568 _1421_ _0294_ _1420_ sg13g2_a21oi_1
Xhold218 _0584_ VPWR VGND net260 sg13g2_dlygate4sd3_1
X_3332_ net271 net569 _1381_ VPWR VGND sg13g2_nor2_1
XFILLER_4_991 VPWR VGND sg13g2_decap_8
Xfanout709 _1963_ net709 VPWR VGND sg13g2_buf_8
X_3263_ VPWR VGND _1279_ _1328_ _1329_ net808 _1330_ _1325_ sg13g2_a221oi_1
X_2214_ VPWR _0516_ _0515_ VGND sg13g2_inv_1
X_3194_ VGND VPWR _1266_ _1267_ _1268_ net578 sg13g2_a21oi_1
XFILLER_38_100 VPWR VGND sg13g2_fill_1
X_2145_ net521 net49 _0448_ VPWR VGND sg13g2_nor2b_2
XFILLER_38_166 VPWR VGND sg13g2_fill_1
X_2076_ VPWR _1955_ net479 VGND sg13g2_inv_1
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_35_873 VPWR VGND sg13g2_fill_2
XFILLER_34_394 VPWR VGND sg13g2_decap_4
XFILLER_14_49 VPWR VGND sg13g2_decap_8
X_2978_ _1123_ _1128_ u_usb_cdc.sie_in_data_ack _1130_ VPWR VGND sg13g2_nand3_1
Xhold730 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\] VPWR VGND
+ net1048 sg13g2_dlygate4sd3_1
XFILLER_2_928 VPWR VGND sg13g2_decap_8
Xhold752 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\] VPWR
+ VGND net1070 sg13g2_dlygate4sd3_1
Xhold741 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[0\] VPWR
+ VGND net1059 sg13g2_dlygate4sd3_1
XFILLER_1_449 VPWR VGND sg13g2_decap_8
XFILLER_29_144 VPWR VGND sg13g2_fill_2
XFILLER_29_155 VPWR VGND sg13g2_fill_2
XFILLER_45_659 VPWR VGND sg13g2_fill_2
XFILLER_38_1012 VPWR VGND sg13g2_decap_8
XFILLER_38_1023 VPWR VGND sg13g2_fill_2
XFILLER_41_832 VPWR VGND sg13g2_fill_1
XFILLER_9_516 VPWR VGND sg13g2_decap_8
XFILLER_41_898 VPWR VGND sg13g2_decap_8
XFILLER_9_527 VPWR VGND sg13g2_fill_1
XFILLER_5_722 VPWR VGND sg13g2_decap_8
XFILLER_5_799 VPWR VGND sg13g2_decap_8
XFILLER_49_921 VPWR VGND sg13g2_decap_8
XFILLER_0_493 VPWR VGND sg13g2_decap_8
XFILLER_49_998 VPWR VGND sg13g2_decap_8
Xhold90 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[42\] VPWR VGND
+ net132 sg13g2_dlygate4sd3_1
XFILLER_36_615 VPWR VGND sg13g2_fill_2
XFILLER_35_147 VPWR VGND sg13g2_decap_8
X_3950_ _1840_ VPWR _1841_ VGND _0585_ _1837_ sg13g2_o21ai_1
X_2901_ net436 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ _1100_ _0115_ VPWR VGND sg13g2_mux2_1
X_3881_ net712 _1737_ _1794_ VPWR VGND sg13g2_nor2_1
X_2832_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net554 _1058_ _0088_ VPWR VGND sg13g2_mux2_1
X_2763_ VGND VPWR net836 _1008_ _1009_ _1006_ sg13g2_a21oi_1
X_2694_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] VPWR _0956_ VGND net622 _2003_ sg13g2_o21ai_1
X_4433_ net696 VGND VPWR net266 u_usb_cdc.u_sie.u_phy_tx.data_q\[3\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_4364_ net695 VGND VPWR _0366_ u_usb_cdc.u_sie.pid_q\[0\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_4295_ net674 VGND VPWR _0297_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[2\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_3315_ net795 net803 net790 _1369_ VPWR VGND sg13g2_a21o_1
X_3246_ net806 net601 _1311_ _1314_ _1315_ VPWR VGND sg13g2_nor4_1
XFILLER_6_1010 VPWR VGND sg13g2_decap_8
X_3177_ _0735_ VPWR _1253_ VGND net768 _1252_ sg13g2_o21ai_1
X_2128_ _2006_ net931 _2004_ VPWR VGND sg13g2_nand2_1
X_2059_ VPWR _1938_ net915 VGND sg13g2_inv_1
XFILLER_25_15 VPWR VGND sg13g2_decap_4
XFILLER_41_139 VPWR VGND sg13g2_fill_2
XFILLER_22_375 VPWR VGND sg13g2_decap_8
XFILLER_41_47 VPWR VGND sg13g2_fill_2
XFILLER_41_36 VPWR VGND sg13g2_fill_2
XFILLER_2_725 VPWR VGND sg13g2_decap_8
Xhold560 u_usb_cdc.bus_reset VPWR VGND net878 sg13g2_dlygate4sd3_1
Xhold571 _0017_ VPWR VGND net889 sg13g2_dlygate4sd3_1
Xhold593 net26 VPWR VGND net911 sg13g2_dlygate4sd3_1
Xhold582 _1723_ VPWR VGND net900 sg13g2_dlygate4sd3_1
XFILLER_46_935 VPWR VGND sg13g2_decap_8
XFILLER_45_456 VPWR VGND sg13g2_fill_2
XFILLER_33_618 VPWR VGND sg13g2_decap_4
XFILLER_25_180 VPWR VGND sg13g2_fill_2
XFILLER_5_541 VPWR VGND sg13g2_fill_2
XFILLER_5_530 VPWR VGND sg13g2_decap_8
X_3100_ _1205_ VPWR _0209_ VGND net708 _1155_ sg13g2_o21ai_1
X_4080_ net654 VGND VPWR net379 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[0\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_49_795 VPWR VGND sg13g2_decap_8
X_3031_ _1164_ net221 _1146_ VPWR VGND sg13g2_nand2_1
XFILLER_36_412 VPWR VGND sg13g2_decap_8
XFILLER_37_968 VPWR VGND sg13g2_decap_8
XFILLER_36_467 VPWR VGND sg13g2_decap_8
X_3933_ _1826_ _2005_ _1824_ VPWR VGND sg13g2_nand2_1
X_3864_ _1739_ VPWR _1783_ VGND net305 _1779_ sg13g2_o21ai_1
X_2815_ _1056_ net542 _1055_ VPWR VGND sg13g2_nand2_2
XFILLER_9_880 VPWR VGND sg13g2_fill_2
X_3795_ _1731_ _1729_ _1730_ VPWR VGND sg13g2_nand2b_1
X_2746_ net423 _0992_ _0993_ VPWR VGND sg13g2_nor2_1
X_2677_ VPWR _0031_ _0944_ VGND sg13g2_inv_1
X_4416_ net729 VGND VPWR _0415_ u_usb_cdc.u_sie.rx_data\[3\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_4347_ net691 VGND VPWR _0349_ u_usb_cdc.sie_out_data\[2\] clknet_leaf_46_clk sg13g2_dfrbpq_2
X_4278_ net693 VGND VPWR net459 u_usb_cdc.u_ctrl_endp.addr_dd\[5\] clknet_leaf_46_clk
+ sg13g2_dfrbpq_1
X_3229_ net817 net321 _1299_ VPWR VGND sg13g2_nor2_1
XFILLER_27_401 VPWR VGND sg13g2_decap_8
XFILLER_14_117 VPWR VGND sg13g2_fill_1
XFILLER_7_839 VPWR VGND sg13g2_fill_1
XFILLER_7_817 VPWR VGND sg13g2_decap_8
XFILLER_2_511 VPWR VGND sg13g2_fill_1
XFILLER_7_2 VPWR VGND sg13g2_fill_1
Xhold390 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[69\] VPWR VGND
+ net432 sg13g2_dlygate4sd3_1
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_42_1019 VPWR VGND sg13g2_decap_8
XFILLER_46_732 VPWR VGND sg13g2_decap_8
XFILLER_19_957 VPWR VGND sg13g2_decap_8
XFILLER_45_231 VPWR VGND sg13g2_fill_1
XFILLER_18_478 VPWR VGND sg13g2_fill_1
XFILLER_34_938 VPWR VGND sg13g2_decap_8
X_2600_ _0874_ _0876_ _0878_ _0880_ _0881_ VPWR VGND sg13g2_nor4_1
X_3580_ net774 _1918_ _1510_ _1554_ _1555_ VPWR VGND sg13g2_nor4_1
X_2531_ net906 VPWR _0826_ VGND _0820_ _0825_ sg13g2_o21ai_1
X_2462_ _0759_ _0758_ _0657_ _0756_ _0688_ VPWR VGND sg13g2_a22oi_1
X_4201_ net662 VGND VPWR net99 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[37\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2393_ net586 net583 net619 _0693_ VPWR VGND sg13g2_nor3_2
XFILLER_3_51 VPWR VGND sg13g2_fill_1
X_4132_ net671 VGND VPWR net127 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[52\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_49_570 VPWR VGND sg13g2_fill_1
X_4063_ net724 VGND VPWR _0034_ u_usb_cdc.u_sie.u_phy_rx.state_q\[2\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_3014_ net823 _1150_ net759 _1153_ VPWR VGND sg13g2_nand3_1
XFILLER_25_938 VPWR VGND sg13g2_fill_2
XFILLER_24_459 VPWR VGND sg13g2_fill_1
XFILLER_33_993 VPWR VGND sg13g2_decap_8
X_3916_ _1810_ u_usb_cdc.u_sie.data_q\[0\] net835 u_usb_cdc.u_sie.pid_q\[0\] net830
+ VPWR VGND sg13g2_a22oi_1
XFILLER_20_610 VPWR VGND sg13g2_decap_8
X_3847_ _1770_ net710 net422 VPWR VGND sg13g2_nand2_1
X_3778_ _1721_ _1720_ net531 net579 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_4_809 VPWR VGND sg13g2_decap_8
X_2729_ VGND VPWR _1902_ _0468_ _0977_ _0466_ sg13g2_a21oi_1
XFILLER_47_529 VPWR VGND sg13g2_fill_2
XFILLER_47_24 VPWR VGND sg13g2_decap_4
XFILLER_27_220 VPWR VGND sg13g2_decap_4
XFILLER_28_776 VPWR VGND sg13g2_fill_1
XFILLER_42_223 VPWR VGND sg13g2_decap_8
XFILLER_27_297 VPWR VGND sg13g2_fill_2
XFILLER_24_982 VPWR VGND sg13g2_decap_8
XFILLER_3_864 VPWR VGND sg13g2_decap_8
XFILLER_2_385 VPWR VGND sg13g2_decap_8
XFILLER_38_529 VPWR VGND sg13g2_decap_8
XFILLER_33_245 VPWR VGND sg13g2_fill_1
XFILLER_18_1021 VPWR VGND sg13g2_decap_8
XFILLER_14_470 VPWR VGND sg13g2_decap_4
XFILLER_30_963 VPWR VGND sg13g2_decap_8
X_3701_ VGND VPWR net794 _1669_ _1670_ net790 sg13g2_a21oi_1
X_3632_ _1604_ net980 net593 VPWR VGND sg13g2_nand2_1
X_3563_ _1538_ _1535_ _1537_ VPWR VGND sg13g2_nand2_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_3494_ _0323_ net573 _1485_ net576 _1946_ VPWR VGND sg13g2_a22oi_1
X_2514_ _1905_ _0734_ _0736_ _0811_ VPWR VGND sg13g2_nor3_1
X_2445_ _0742_ net953 _0692_ VPWR VGND sg13g2_nand2_1
X_4115_ net657 VGND VPWR net455 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[35\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2376_ _0676_ net736 _0675_ VPWR VGND sg13g2_nand2_1
XFILLER_29_507 VPWR VGND sg13g2_decap_4
X_4046_ net694 VGND VPWR net414 u_usb_cdc.u_sie.phy_state_q\[2\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_37_540 VPWR VGND sg13g2_fill_2
XFILLER_40_727 VPWR VGND sg13g2_decap_8
XFILLER_40_749 VPWR VGND sg13g2_fill_1
XFILLER_0_801 VPWR VGND sg13g2_decap_8
XFILLER_48_805 VPWR VGND sg13g2_decap_8
XFILLER_0_878 VPWR VGND sg13g2_decap_8
XFILLER_43_587 VPWR VGND sg13g2_decap_4
XFILLER_12_930 VPWR VGND sg13g2_decap_8
XFILLER_8_945 VPWR VGND sg13g2_decap_8
XFILLER_3_661 VPWR VGND sg13g2_decap_8
X_2230_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] u_usb_cdc.u_ctrl_endp.max_length_q\[6\]
+ _0532_ VPWR VGND sg13g2_xor2_1
X_2161_ _0463_ net755 u_usb_cdc.addr\[3\] VPWR VGND sg13g2_xnor2_1
XFILLER_17_4 VPWR VGND sg13g2_fill_2
X_2092_ VPWR _1970_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[43\]
+ VGND sg13g2_inv_1
XFILLER_22_727 VPWR VGND sg13g2_fill_1
X_2994_ _1140_ net82 net614 VPWR VGND sg13g2_nand2_1
X_3615_ VGND VPWR net791 _1587_ _1588_ _1913_ sg13g2_a21oi_1
X_3546_ _1513_ _1518_ _1509_ _1522_ VPWR VGND _1521_ sg13g2_nand4_1
X_3477_ _1473_ net289 net594 VPWR VGND sg13g2_nand2_1
X_2428_ _0726_ net937 VPWR VGND net346 sg13g2_nand2b_2
X_2359_ net586 net583 net620 _0659_ VPWR VGND sg13g2_nor3_1
XFILLER_29_315 VPWR VGND sg13g2_fill_2
X_4029_ net665 VGND VPWR net950 u_usb_cdc.u_ctrl_endp.req_q\[9\] clknet_leaf_49_clk
+ sg13g2_dfrbpq_1
XFILLER_25_543 VPWR VGND sg13g2_fill_1
XFILLER_37_381 VPWR VGND sg13g2_fill_1
XFILLER_44_69 VPWR VGND sg13g2_fill_1
XFILLER_40_524 VPWR VGND sg13g2_fill_2
XFILLER_12_237 VPWR VGND sg13g2_fill_1
XFILLER_40_546 VPWR VGND sg13g2_decap_8
XFILLER_21_760 VPWR VGND sg13g2_decap_4
XFILLER_5_904 VPWR VGND sg13g2_decap_8
XFILLER_4_458 VPWR VGND sg13g2_decap_8
XFILLER_0_675 VPWR VGND sg13g2_decap_8
XFILLER_44_885 VPWR VGND sg13g2_decap_8
XFILLER_43_351 VPWR VGND sg13g2_fill_2
XFILLER_16_576 VPWR VGND sg13g2_fill_2
XFILLER_8_731 VPWR VGND sg13g2_decap_8
XFILLER_8_742 VPWR VGND sg13g2_fill_1
XFILLER_12_793 VPWR VGND sg13g2_fill_2
XFILLER_7_274 VPWR VGND sg13g2_decap_8
Xhold208 u_usb_cdc.u_sie.addr_q\[6\] VPWR VGND net250 sg13g2_dlygate4sd3_1
X_4380_ net722 VGND VPWR net332 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[1\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_2
X_3400_ u_usb_cdc.sie_out_data\[6\] _1408_ _1421_ VPWR VGND sg13g2_nor2_1
Xhold219 _0596_ VPWR VGND net261 sg13g2_dlygate4sd3_1
XFILLER_4_970 VPWR VGND sg13g2_decap_8
X_3331_ VGND VPWR net718 net569 _0265_ _1380_ sg13g2_a21oi_1
X_3262_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[5\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[13\]
+ net818 _1329_ VPWR VGND sg13g2_mux2_1
X_2213_ _0515_ _1946_ _0512_ VPWR VGND sg13g2_xnor2_1
X_3193_ _1267_ _0606_ _1265_ net983 net749 VPWR VGND sg13g2_a22oi_1
XFILLER_39_613 VPWR VGND sg13g2_fill_1
X_2144_ net360 _1934_ _0445_ _0446_ _0447_ VPWR VGND sg13g2_and4_1
XFILLER_39_668 VPWR VGND sg13g2_decap_4
X_2075_ VPWR _1954_ u_usb_cdc.addr\[0\] VGND sg13g2_inv_1
XFILLER_14_28 VPWR VGND sg13g2_fill_1
X_2977_ _1129_ net1034 _1128_ VPWR VGND sg13g2_nand2_1
XFILLER_2_907 VPWR VGND sg13g2_decap_8
Xhold720 _0855_ VPWR VGND net1038 sg13g2_dlygate4sd3_1
Xhold731 u_usb_cdc.clk_gate_q VPWR VGND net1049 sg13g2_dlygate4sd3_1
Xhold742 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[2\] VPWR VGND net1060 sg13g2_dlygate4sd3_1
XFILLER_1_428 VPWR VGND sg13g2_decap_8
X_3529_ VGND VPWR net780 _0651_ _1505_ net776 sg13g2_a21oi_1
XFILLER_39_25 VPWR VGND sg13g2_fill_2
XFILLER_44_126 VPWR VGND sg13g2_decap_4
XFILLER_29_189 VPWR VGND sg13g2_fill_1
XFILLER_25_395 VPWR VGND sg13g2_fill_1
XFILLER_40_376 VPWR VGND sg13g2_fill_1
XFILLER_5_701 VPWR VGND sg13g2_decap_8
XFILLER_5_778 VPWR VGND sg13g2_decap_8
XFILLER_45_1017 VPWR VGND sg13g2_decap_8
XFILLER_49_900 VPWR VGND sg13g2_decap_8
XFILLER_45_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_472 VPWR VGND sg13g2_decap_8
XFILLER_1_995 VPWR VGND sg13g2_decap_8
XFILLER_49_977 VPWR VGND sg13g2_decap_8
Xhold80 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[10\] VPWR VGND
+ net122 sg13g2_dlygate4sd3_1
Xhold91 _0209_ VPWR VGND net133 sg13g2_dlygate4sd3_1
XFILLER_35_137 VPWR VGND sg13g2_fill_1
X_2900_ net828 net827 net615 _1100_ VPWR VGND sg13g2_nor3_2
X_3880_ VGND VPWR net52 _1791_ _0401_ _1793_ sg13g2_a21oi_1
XFILLER_31_387 VPWR VGND sg13g2_fill_2
X_2831_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net397 _1058_ _0087_ VPWR VGND sg13g2_mux2_1
X_2762_ _1008_ _1004_ _1007_ VPWR VGND sg13g2_nand2_1
X_4432_ net696 VGND VPWR net212 u_usb_cdc.u_sie.u_phy_tx.data_q\[2\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_2693_ _0953_ net702 net557 _0036_ VPWR VGND sg13g2_nor3_1
X_4363_ net641 VGND VPWR net934 net28 clknet_leaf_11_clk sg13g2_dfrbpq_2
X_4294_ net674 VGND VPWR _0296_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[1\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
X_3314_ net795 net790 net803 _1368_ VPWR VGND sg13g2_nand3_1
X_3245_ VPWR VGND _1309_ net807 _1313_ net809 _1314_ _1312_ sg13g2_a221oi_1
X_3176_ _1241_ _1247_ _1251_ _1252_ VPWR VGND sg13g2_nor3_1
XFILLER_27_605 VPWR VGND sg13g2_fill_1
XFILLER_27_627 VPWR VGND sg13g2_decap_4
XFILLER_39_454 VPWR VGND sg13g2_fill_1
X_2127_ _2005_ _1994_ net705 VPWR VGND sg13g2_nand2_1
XFILLER_27_638 VPWR VGND sg13g2_decap_4
X_2058_ _1937_ net935 VPWR VGND sg13g2_inv_2
XFILLER_35_693 VPWR VGND sg13g2_fill_2
XFILLER_10_527 VPWR VGND sg13g2_fill_1
XFILLER_2_704 VPWR VGND sg13g2_decap_8
Xhold550 u_usb_cdc.u_ctrl_endp.req_q\[1\] VPWR VGND net868 sg13g2_dlygate4sd3_1
Xhold572 u_usb_cdc.u_ctrl_endp.max_length_q\[6\] VPWR VGND net890 sg13g2_dlygate4sd3_1
Xhold561 _0402_ VPWR VGND net879 sg13g2_dlygate4sd3_1
Xhold583 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\] VPWR VGND
+ net901 sg13g2_dlygate4sd3_1
Xhold594 _0363_ VPWR VGND net912 sg13g2_dlygate4sd3_1
XFILLER_49_218 VPWR VGND sg13g2_fill_1
XFILLER_1_269 VPWR VGND sg13g2_fill_1
XFILLER_46_914 VPWR VGND sg13g2_decap_8
XFILLER_18_616 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_52_clk clknet_3_1__leaf_clk clknet_leaf_52_clk VPWR VGND sg13g2_buf_8
XFILLER_13_354 VPWR VGND sg13g2_decap_4
XFILLER_14_877 VPWR VGND sg13g2_fill_2
XFILLER_1_792 VPWR VGND sg13g2_decap_8
XFILLER_49_774 VPWR VGND sg13g2_decap_8
X_3030_ _1162_ VPWR _0181_ VGND net821 _1163_ sg13g2_o21ai_1
XFILLER_37_947 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_43_clk clknet_3_4__leaf_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
X_3932_ net623 VPWR _1825_ VGND _1993_ _1034_ sg13g2_o21ai_1
X_3863_ net305 _1779_ _1782_ VPWR VGND sg13g2_and2_1
XFILLER_20_825 VPWR VGND sg13g2_fill_1
XFILLER_32_652 VPWR VGND sg13g2_decap_8
X_2814_ VGND VPWR _1055_ _1054_ net714 sg13g2_or2_1
X_3794_ _0936_ VPWR _1730_ VGND _0441_ _0915_ sg13g2_o21ai_1
XFILLER_8_380 VPWR VGND sg13g2_fill_2
X_2745_ _0992_ net518 _0991_ VPWR VGND sg13g2_nand2_1
XFILLER_9_892 VPWR VGND sg13g2_fill_2
X_2676_ _0944_ net635 _0943_ net704 net515 VPWR VGND sg13g2_a22oi_1
X_4415_ net729 VGND VPWR _0414_ u_usb_cdc.u_sie.rx_data\[2\] clknet_leaf_34_clk sg13g2_dfrbpq_2
X_4346_ net682 VGND VPWR _0348_ u_usb_cdc.sie_out_data\[1\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_28_1012 VPWR VGND sg13g2_decap_8
X_4277_ net693 VGND VPWR net385 u_usb_cdc.u_ctrl_endp.addr_dd\[4\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_3228_ net817 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[34\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[42\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[50\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[58\] net811 _1298_
+ VPWR VGND sg13g2_mux4_1
XFILLER_28_914 VPWR VGND sg13g2_decap_8
X_3159_ _1237_ net116 _1230_ VPWR VGND sg13g2_nand2_1
XFILLER_42_405 VPWR VGND sg13g2_fill_2
XFILLER_23_641 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_34_clk clknet_3_7__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
XFILLER_22_151 VPWR VGND sg13g2_decap_4
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_22_162 VPWR VGND sg13g2_decap_8
XFILLER_10_357 VPWR VGND sg13g2_decap_8
XFILLER_2_523 VPWR VGND sg13g2_fill_2
Xhold380 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[11\] VPWR VGND net422 sg13g2_dlygate4sd3_1
XFILLER_2_578 VPWR VGND sg13g2_decap_8
Xhold391 _0152_ VPWR VGND net433 sg13g2_dlygate4sd3_1
XFILLER_46_711 VPWR VGND sg13g2_decap_8
XFILLER_46_788 VPWR VGND sg13g2_decap_8
XFILLER_14_641 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_25_clk clknet_3_6__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
X_2530_ _0822_ _0823_ _0821_ _0825_ VPWR VGND _0824_ sg13g2_nand4_1
XFILLER_6_884 VPWR VGND sg13g2_decap_8
X_2461_ _0758_ _0751_ _0752_ VPWR VGND sg13g2_nand2_1
X_4200_ net664 VGND VPWR net241 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[36\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_2392_ _0678_ _0691_ _0663_ _0692_ VPWR VGND sg13g2_nand3_1
X_4131_ net651 VGND VPWR net160 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[51\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_4062_ net724 VGND VPWR net344 u_usb_cdc.u_sie.u_phy_rx.state_q\[1\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_2
X_3013_ _1152_ net216 _1146_ VPWR VGND sg13g2_nand2_1
XFILLER_3_1025 VPWR VGND sg13g2_decap_4
XFILLER_37_711 VPWR VGND sg13g2_decap_4
XFILLER_37_777 VPWR VGND sg13g2_fill_1
XFILLER_24_405 VPWR VGND sg13g2_fill_2
XFILLER_36_254 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_16_clk clknet_3_2__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_3915_ _1809_ _1952_ net831 _1938_ net838 VPWR VGND sg13g2_a22oi_1
XFILLER_33_972 VPWR VGND sg13g2_decap_8
X_3846_ _1767_ VPWR _0391_ VGND _1768_ _1769_ sg13g2_o21ai_1
XFILLER_20_655 VPWR VGND sg13g2_fill_2
X_3777_ _1718_ _1719_ _1720_ VPWR VGND sg13g2_nor2b_2
X_2728_ _0976_ _0601_ _0469_ VPWR VGND sg13g2_nand2b_1
X_2659_ net618 _0726_ u_usb_cdc.u_ctrl_endp.in_dir_q _0929_ VPWR VGND sg13g2_nand3_1
X_4329_ net695 VGND VPWR _0331_ u_usb_cdc.u_sie.crc16_q\[8\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_47_508 VPWR VGND sg13g2_decap_8
XFILLER_47_47 VPWR VGND sg13g2_fill_2
XFILLER_16_917 VPWR VGND sg13g2_fill_2
XFILLER_43_725 VPWR VGND sg13g2_fill_1
XFILLER_15_416 VPWR VGND sg13g2_fill_1
XFILLER_15_427 VPWR VGND sg13g2_fill_2
XFILLER_28_799 VPWR VGND sg13g2_decap_4
XFILLER_23_471 VPWR VGND sg13g2_decap_8
XFILLER_23_482 VPWR VGND sg13g2_decap_4
XFILLER_23_493 VPWR VGND sg13g2_fill_1
XFILLER_10_132 VPWR VGND sg13g2_decap_4
XFILLER_10_176 VPWR VGND sg13g2_decap_4
XFILLER_12_83 VPWR VGND sg13g2_fill_2
XFILLER_3_843 VPWR VGND sg13g2_decap_8
XFILLER_2_364 VPWR VGND sg13g2_decap_8
Xfanout690 net701 net690 VPWR VGND sg13g2_buf_8
XFILLER_22_909 VPWR VGND sg13g2_fill_1
XFILLER_33_224 VPWR VGND sg13g2_fill_2
XFILLER_34_736 VPWR VGND sg13g2_decap_4
XFILLER_18_1000 VPWR VGND sg13g2_decap_8
XFILLER_30_920 VPWR VGND sg13g2_fill_2
X_3700_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[23\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[31\]
+ net801 _1669_ VPWR VGND sg13g2_mux2_1
X_3631_ _1582_ VPWR _0342_ VGND _1602_ _1603_ sg13g2_o21ai_1
X_3562_ VGND VPWR net792 _1536_ _1537_ _1913_ sg13g2_a21oi_1
X_2513_ _1930_ _0699_ _0743_ _0810_ VPWR VGND sg13g2_nor3_1
X_3493_ _0514_ _0500_ _1485_ VPWR VGND sg13g2_xor2_1
X_2444_ _0725_ VPWR _0005_ VGND _0732_ _0741_ sg13g2_o21ai_1
Xclkbuf_leaf_5_clk clknet_3_0__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_2375_ net787 net715 _0655_ _0675_ VPWR VGND sg13g2_nor3_2
X_4114_ net656 VGND VPWR net447 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[34\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_25_1026 VPWR VGND sg13g2_fill_2
X_4045_ net694 VGND VPWR net1051 u_usb_cdc.u_sie.phy_state_q\[1\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
XFILLER_37_552 VPWR VGND sg13g2_fill_1
XFILLER_25_703 VPWR VGND sg13g2_fill_1
XFILLER_37_585 VPWR VGND sg13g2_decap_4
XFILLER_40_706 VPWR VGND sg13g2_decap_8
XFILLER_20_441 VPWR VGND sg13g2_fill_1
X_3829_ VGND VPWR net600 _1753_ _1757_ net172 sg13g2_a21oi_1
XFILLER_20_485 VPWR VGND sg13g2_fill_2
XFILLER_4_618 VPWR VGND sg13g2_fill_1
XFILLER_0_857 VPWR VGND sg13g2_decap_8
XFILLER_47_349 VPWR VGND sg13g2_fill_2
XFILLER_15_213 VPWR VGND sg13g2_fill_1
XFILLER_28_596 VPWR VGND sg13g2_decap_4
XFILLER_43_577 VPWR VGND sg13g2_fill_1
XFILLER_8_924 VPWR VGND sg13g2_decap_8
XFILLER_12_986 VPWR VGND sg13g2_decap_8
XFILLER_48_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_640 VPWR VGND sg13g2_decap_8
X_2160_ u_usb_cdc.addr\[0\] net760 _0462_ VPWR VGND sg13g2_xor2_1
X_2091_ VPWR _1969_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[42\]
+ VGND sg13g2_inv_1
XFILLER_38_349 VPWR VGND sg13g2_fill_2
XFILLER_46_360 VPWR VGND sg13g2_fill_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
X_2993_ _1139_ VPWR _0168_ VGND net720 net613 sg13g2_o21ai_1
X_3614_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[51\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[59\]
+ net798 _1587_ VPWR VGND sg13g2_mux2_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
X_3545_ _0552_ VPWR _1521_ VGND _1519_ _1520_ sg13g2_o21ai_1
X_3476_ VGND VPWR _1921_ _1471_ _0318_ _1468_ sg13g2_a21oi_1
X_2427_ net971 VPWR _0725_ VGND _0720_ _0721_ sg13g2_o21ai_1
X_2358_ _0658_ u_usb_cdc.u_ctrl_endp.state_q\[2\] _0605_ VPWR VGND sg13g2_nand2_1
X_2289_ _0591_ _1904_ net743 VPWR VGND sg13g2_nand2_1
X_4028_ net666 VGND VPWR net846 u_usb_cdc.u_ctrl_endp.req_q\[8\] clknet_leaf_49_clk
+ sg13g2_dfrbpq_2
XFILLER_25_522 VPWR VGND sg13g2_fill_1
XFILLER_25_588 VPWR VGND sg13g2_fill_2
XFILLER_20_293 VPWR VGND sg13g2_fill_1
XFILLER_0_654 VPWR VGND sg13g2_decap_8
XFILLER_48_625 VPWR VGND sg13g2_fill_2
XFILLER_44_864 VPWR VGND sg13g2_decap_8
XFILLER_16_599 VPWR VGND sg13g2_decap_8
XFILLER_31_514 VPWR VGND sg13g2_decap_8
XFILLER_12_783 VPWR VGND sg13g2_fill_2
XFILLER_8_776 VPWR VGND sg13g2_decap_8
Xhold209 _0312_ VPWR VGND net251 sg13g2_dlygate4sd3_1
X_3330_ net341 net569 _1380_ VPWR VGND sg13g2_nor2_1
XFILLER_3_470 VPWR VGND sg13g2_fill_1
X_3261_ _1278_ _1326_ _1327_ _1328_ VPWR VGND sg13g2_nor3_1
X_2212_ _0514_ _0508_ _0513_ VPWR VGND sg13g2_xnor2_1
X_3192_ _1266_ _0735_ _1245_ VPWR VGND sg13g2_nand2_1
XFILLER_22_1018 VPWR VGND sg13g2_decap_8
X_2143_ net428 net527 _0446_ VPWR VGND sg13g2_nor2_1
XFILLER_38_135 VPWR VGND sg13g2_decap_4
XFILLER_39_658 VPWR VGND sg13g2_fill_2
XFILLER_38_157 VPWR VGND sg13g2_decap_8
X_2074_ _1953_ net349 VPWR VGND sg13g2_inv_2
XFILLER_19_371 VPWR VGND sg13g2_decap_4
XFILLER_34_341 VPWR VGND sg13g2_fill_1
X_2976_ _1128_ u_usb_cdc.sie_in_req net631 VPWR VGND sg13g2_nand2_2
Xhold721 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ VPWR VGND net1039 sg13g2_dlygate4sd3_1
Xhold710 _0260_ VPWR VGND net1028 sg13g2_dlygate4sd3_1
XFILLER_1_407 VPWR VGND sg13g2_decap_8
Xhold732 u_usb_cdc.u_sie.phy_state_q\[1\] VPWR VGND net1050 sg13g2_dlygate4sd3_1
Xhold743 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[3\] VPWR VGND net1061 sg13g2_dlygate4sd3_1
X_3528_ _1504_ net780 _0651_ VPWR VGND sg13g2_nand2_1
X_3459_ _1460_ net937 _1456_ _0313_ VPWR VGND sg13g2_mux2_1
XFILLER_45_617 VPWR VGND sg13g2_fill_2
XFILLER_29_179 VPWR VGND sg13g2_fill_1
XFILLER_26_831 VPWR VGND sg13g2_decap_4
XFILLER_26_897 VPWR VGND sg13g2_fill_2
XFILLER_40_355 VPWR VGND sg13g2_decap_8
XFILLER_5_757 VPWR VGND sg13g2_decap_8
XFILLER_0_451 VPWR VGND sg13g2_decap_8
XFILLER_1_974 VPWR VGND sg13g2_decap_8
XFILLER_49_956 VPWR VGND sg13g2_decap_8
Xhold81 _0177_ VPWR VGND net123 sg13g2_dlygate4sd3_1
Xhold92 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[69\] VPWR VGND
+ net134 sg13g2_dlygate4sd3_1
Xhold70 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[47\] VPWR VGND
+ net112 sg13g2_dlygate4sd3_1
XFILLER_48_488 VPWR VGND sg13g2_decap_8
XFILLER_29_691 VPWR VGND sg13g2_fill_1
XFILLER_36_639 VPWR VGND sg13g2_fill_2
XFILLER_16_341 VPWR VGND sg13g2_decap_8
X_2830_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net407 _1058_ _0086_ VPWR VGND sg13g2_mux2_1
XFILLER_32_856 VPWR VGND sg13g2_fill_2
XFILLER_12_591 VPWR VGND sg13g2_fill_1
X_2761_ net762 net1011 _1989_ _0882_ _1007_ VPWR VGND sg13g2_nor4_1
X_2692_ VGND VPWR net623 net705 _0955_ net556 sg13g2_a21oi_1
X_4431_ net698 VGND VPWR _0422_ u_usb_cdc.u_sie.u_phy_tx.data_q\[1\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_4362_ net641 VGND VPWR net963 net27 clknet_leaf_11_clk sg13g2_dfrbpq_2
X_4293_ net674 VGND VPWR _0295_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[0\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
X_3313_ net1027 VPWR _0260_ VGND _1358_ _1366_ sg13g2_o21ai_1
X_3244_ VGND VPWR net813 _1978_ _1313_ net809 sg13g2_a21oi_1
XFILLER_20_0 VPWR VGND sg13g2_fill_1
X_3175_ _1250_ net806 _1251_ VPWR VGND sg13g2_xor2_1
XFILLER_26_105 VPWR VGND sg13g2_fill_2
XFILLER_26_127 VPWR VGND sg13g2_decap_8
X_2126_ _1993_ _2003_ _2004_ VPWR VGND sg13g2_nor2_1
X_2057_ VPWR _1936_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] VGND sg13g2_inv_1
XFILLER_25_28 VPWR VGND sg13g2_fill_1
XFILLER_22_322 VPWR VGND sg13g2_fill_1
XFILLER_22_355 VPWR VGND sg13g2_decap_8
X_2959_ net432 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ _1121_ _0152_ VPWR VGND sg13g2_mux2_1
XFILLER_41_49 VPWR VGND sg13g2_fill_1
Xhold551 _0002_ VPWR VGND net869 sg13g2_dlygate4sd3_1
Xhold562 u_usb_cdc.addr\[1\] VPWR VGND net880 sg13g2_dlygate4sd3_1
Xhold540 net18 VPWR VGND net858 sg13g2_dlygate4sd3_1
Xhold584 _0157_ VPWR VGND net902 sg13g2_dlygate4sd3_1
Xhold573 _0294_ VPWR VGND net891 sg13g2_dlygate4sd3_1
Xhold595 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\] VPWR VGND net913 sg13g2_dlygate4sd3_1
XFILLER_25_182 VPWR VGND sg13g2_fill_1
XFILLER_41_675 VPWR VGND sg13g2_decap_8
XFILLER_41_653 VPWR VGND sg13g2_fill_1
XFILLER_13_377 VPWR VGND sg13g2_fill_1
XFILLER_14_889 VPWR VGND sg13g2_decap_8
XFILLER_40_163 VPWR VGND sg13g2_fill_2
XFILLER_1_771 VPWR VGND sg13g2_decap_8
XFILLER_49_753 VPWR VGND sg13g2_decap_8
XFILLER_37_926 VPWR VGND sg13g2_decap_8
XFILLER_36_447 VPWR VGND sg13g2_decap_8
X_3931_ VGND VPWR _1999_ _1824_ _1033_ net702 sg13g2_a21oi_2
X_3862_ _1781_ net711 net305 VPWR VGND sg13g2_nand2_1
XFILLER_31_130 VPWR VGND sg13g2_fill_2
XFILLER_31_163 VPWR VGND sg13g2_fill_2
XFILLER_32_697 VPWR VGND sg13g2_fill_2
X_2813_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq
+ VPWR _1054_ VGND _1051_ _1053_ sg13g2_o21ai_1
X_3793_ _0441_ VPWR _1729_ VGND _0918_ _1728_ sg13g2_o21ai_1
X_2744_ net341 net271 _0991_ VPWR VGND sg13g2_nor2_1
X_2675_ _0942_ VPWR _0943_ VGND net351 _0455_ sg13g2_o21ai_1
X_4414_ net729 VGND VPWR _0413_ u_usb_cdc.u_sie.rx_data\[1\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_4345_ net681 VGND VPWR _0347_ u_usb_cdc.sie_out_data\[0\] clknet_leaf_46_clk sg13g2_dfrbpq_2
X_4276_ net679 VGND VPWR _0278_ u_usb_cdc.u_ctrl_endp.addr_dd\[3\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
X_3227_ _0244_ _1297_ _1295_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_904 VPWR VGND sg13g2_decap_4
XFILLER_39_230 VPWR VGND sg13g2_fill_1
X_3158_ _1236_ VPWR _0236_ VGND _1178_ _1229_ sg13g2_o21ai_1
XFILLER_36_16 VPWR VGND sg13g2_decap_4
X_2109_ net767 u_usb_cdc.endp\[2\] _1987_ VPWR VGND sg13g2_nor2_1
XFILLER_27_458 VPWR VGND sg13g2_decap_8
XFILLER_43_929 VPWR VGND sg13g2_decap_8
X_3089_ _1199_ VPWR _0204_ VGND _1898_ net607 sg13g2_o21ai_1
XFILLER_35_1006 VPWR VGND sg13g2_decap_8
XFILLER_10_336 VPWR VGND sg13g2_decap_4
XFILLER_2_502 VPWR VGND sg13g2_fill_2
Xhold381 u_usb_cdc.u_ctrl_endp.endp_q\[1\] VPWR VGND net423 sg13g2_dlygate4sd3_1
XFILLER_2_557 VPWR VGND sg13g2_decap_8
Xhold370 net14 VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold392 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[57\] VPWR VGND
+ net434 sg13g2_dlygate4sd3_1
XFILLER_18_414 VPWR VGND sg13g2_fill_1
XFILLER_46_767 VPWR VGND sg13g2_decap_8
XFILLER_42_984 VPWR VGND sg13g2_decap_8
XFILLER_41_494 VPWR VGND sg13g2_decap_8
XFILLER_13_174 VPWR VGND sg13g2_decap_8
XFILLER_9_167 VPWR VGND sg13g2_fill_1
XFILLER_6_863 VPWR VGND sg13g2_decap_8
X_2460_ VGND VPWR _0673_ _0685_ _0757_ _0751_ sg13g2_a21oi_1
XFILLER_5_395 VPWR VGND sg13g2_decap_8
X_4130_ net650 VGND VPWR net125 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[50\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2391_ _0679_ _0684_ _0687_ _0690_ _0691_ VPWR VGND sg13g2_nor4_1
XFILLER_49_561 VPWR VGND sg13g2_decap_8
X_4061_ net724 VGND VPWR _0065_ _0052_ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3012_ _1147_ VPWR _0175_ VGND net821 _1151_ sg13g2_o21ai_1
XFILLER_3_1004 VPWR VGND sg13g2_decap_8
XFILLER_33_951 VPWR VGND sg13g2_decap_8
X_3914_ net748 net702 _1808_ VPWR VGND sg13g2_nor2_1
X_3845_ net600 VPWR _1769_ VGND net303 _1765_ sg13g2_o21ai_1
X_3776_ _1937_ _0933_ _1719_ VPWR VGND sg13g2_nor2_1
X_2727_ u_usb_cdc.bus_reset net722 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.rstn VPWR
+ VGND sg13g2_nor2b_1
X_2658_ net868 VPWR _0928_ VGND _0840_ _0927_ sg13g2_o21ai_1
X_2589_ _0868_ VPWR _0020_ VGND _0469_ net582 sg13g2_o21ai_1
X_4328_ net688 VGND VPWR net883 u_usb_cdc.u_sie.crc16_q\[7\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_4259_ net683 VGND VPWR net990 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[2\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_41_1010 VPWR VGND sg13g2_decap_8
XFILLER_6_104 VPWR VGND sg13g2_fill_2
XFILLER_11_689 VPWR VGND sg13g2_fill_2
XFILLER_3_822 VPWR VGND sg13g2_decap_8
XFILLER_3_899 VPWR VGND sg13g2_decap_8
Xfanout680 net682 net680 VPWR VGND sg13g2_buf_2
Xfanout691 net700 net691 VPWR VGND sg13g2_buf_8
XFILLER_46_542 VPWR VGND sg13g2_fill_2
XFILLER_34_759 VPWR VGND sg13g2_decap_8
XFILLER_14_450 VPWR VGND sg13g2_decap_8
XFILLER_30_998 VPWR VGND sg13g2_decap_8
X_3630_ net597 VPWR _1603_ VGND net966 net624 sg13g2_o21ai_1
X_3561_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[49\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[57\]
+ net797 _1536_ VPWR VGND sg13g2_mux2_1
X_2512_ VGND VPWR _0695_ _0787_ _0809_ _0808_ sg13g2_a21oi_1
XFILLER_5_181 VPWR VGND sg13g2_fill_1
X_3492_ net840 net836 net577 _1484_ VPWR VGND sg13g2_nor3_2
X_2443_ _0741_ _0740_ VPWR VGND _0737_ sg13g2_nand2b_2
X_2374_ VPWR _0674_ _0673_ VGND sg13g2_inv_1
XFILLER_25_1005 VPWR VGND sg13g2_decap_8
X_4113_ net653 VGND VPWR net472 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[33\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4044_ net694 VGND VPWR net262 _0050_ clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_21_932 VPWR VGND sg13g2_fill_2
XFILLER_21_954 VPWR VGND sg13g2_fill_1
X_3828_ VGND VPWR _1981_ _1756_ _0386_ _1755_ sg13g2_a21oi_1
X_3759_ _1702_ _1704_ _1701_ _1705_ VPWR VGND sg13g2_nand3_1
XFILLER_0_836 VPWR VGND sg13g2_decap_8
XFILLER_28_531 VPWR VGND sg13g2_fill_2
XFILLER_16_715 VPWR VGND sg13g2_fill_2
XFILLER_8_903 VPWR VGND sg13g2_decap_8
XFILLER_11_420 VPWR VGND sg13g2_fill_1
XFILLER_12_965 VPWR VGND sg13g2_decap_8
XFILLER_7_402 VPWR VGND sg13g2_fill_2
XFILLER_3_696 VPWR VGND sg13g2_decap_8
XFILLER_39_818 VPWR VGND sg13g2_fill_1
XFILLER_17_6 VPWR VGND sg13g2_fill_1
X_2090_ VPWR _1968_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[41\]
+ VGND sg13g2_inv_1
XFILLER_47_884 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_1018 VPWR VGND sg13g2_decap_8
XFILLER_46_394 VPWR VGND sg13g2_decap_4
X_2992_ _1139_ net97 net613 VPWR VGND sg13g2_nand2_1
XFILLER_9_63 VPWR VGND sg13g2_fill_2
X_3613_ _1585_ VPWR _1586_ VGND net800 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[35\]
+ sg13g2_o21ai_1
X_3544_ VGND VPWR net787 net716 _1520_ _0543_ sg13g2_a21oi_1
X_3475_ _1468_ net508 _1472_ _0317_ VPWR VGND sg13g2_nor3_1
X_2426_ _0724_ net738 _0723_ VPWR VGND sg13g2_nand2_2
X_2357_ _0649_ _0652_ _0657_ VPWR VGND sg13g2_nor2_1
X_2288_ _0589_ VPWR _0590_ VGND _0585_ _0587_ sg13g2_o21ai_1
X_4027_ net676 VGND VPWR net922 u_usb_cdc.u_ctrl_endp.req_q\[7\] clknet_leaf_50_clk
+ sg13g2_dfrbpq_2
XFILLER_25_501 VPWR VGND sg13g2_decap_4
XFILLER_38_862 VPWR VGND sg13g2_fill_2
XFILLER_38_884 VPWR VGND sg13g2_decap_8
XFILLER_12_217 VPWR VGND sg13g2_fill_2
XFILLER_5_939 VPWR VGND sg13g2_decap_8
XFILLER_0_633 VPWR VGND sg13g2_decap_8
XFILLER_44_843 VPWR VGND sg13g2_decap_8
XFILLER_43_353 VPWR VGND sg13g2_fill_1
XFILLER_16_545 VPWR VGND sg13g2_decap_8
XFILLER_16_578 VPWR VGND sg13g2_fill_1
XFILLER_15_1026 VPWR VGND sg13g2_fill_2
XFILLER_8_755 VPWR VGND sg13g2_decap_8
X_3260_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[29\] net818
+ _1327_ VPWR VGND sg13g2_nor2b_1
X_2211_ _0513_ _0509_ _0512_ VPWR VGND sg13g2_xnor2_1
X_3191_ _1264_ VPWR _1265_ VGND net768 net709 sg13g2_o21ai_1
XFILLER_39_626 VPWR VGND sg13g2_decap_4
X_2142_ _1935_ net899 net862 net908 _0445_ VPWR VGND sg13g2_nor4_1
X_2073_ _1952_ net882 VPWR VGND sg13g2_inv_2
XFILLER_35_821 VPWR VGND sg13g2_fill_1
X_2975_ _1052_ net1020 _1055_ _0162_ VPWR VGND sg13g2_mux2_1
XFILLER_30_581 VPWR VGND sg13g2_decap_8
XFILLER_30_592 VPWR VGND sg13g2_fill_1
Xhold711 u_usb_cdc.u_ctrl_endp.req_q\[5\] VPWR VGND net1029 sg13g2_dlygate4sd3_1
Xhold700 u_usb_cdc.u_sie.pid_q\[3\] VPWR VGND net1018 sg13g2_dlygate4sd3_1
Xhold744 u_usb_cdc.sie_out_data\[2\] VPWR VGND net1062 sg13g2_dlygate4sd3_1
Xhold733 _0020_ VPWR VGND net1051 sg13g2_dlygate4sd3_1
Xhold722 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ VPWR VGND net1040 sg13g2_dlygate4sd3_1
X_3527_ _1503_ net770 net773 VPWR VGND sg13g2_nand2b_1
X_3458_ _1459_ VPWR _1460_ VGND net415 _1932_ sg13g2_o21ai_1
XFILLER_39_27 VPWR VGND sg13g2_fill_1
X_2409_ net753 net754 net751 _0707_ VGND VPWR net752 sg13g2_nor4_2
X_3389_ VGND VPWR net567 _1413_ _0290_ _1412_ sg13g2_a21oi_1
XFILLER_29_125 VPWR VGND sg13g2_decap_4
XFILLER_13_537 VPWR VGND sg13g2_decap_8
XFILLER_25_386 VPWR VGND sg13g2_decap_8
XFILLER_5_736 VPWR VGND sg13g2_decap_8
XFILLER_20_84 VPWR VGND sg13g2_fill_1
XFILLER_0_430 VPWR VGND sg13g2_decap_8
XFILLER_1_953 VPWR VGND sg13g2_decap_8
XFILLER_49_935 VPWR VGND sg13g2_decap_8
Xhold82 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[50\] VPWR VGND
+ net124 sg13g2_dlygate4sd3_1
Xhold60 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[11\] VPWR VGND
+ net102 sg13g2_dlygate4sd3_1
Xhold71 _0214_ VPWR VGND net113 sg13g2_dlygate4sd3_1
Xhold93 _0236_ VPWR VGND net135 sg13g2_dlygate4sd3_1
XFILLER_43_172 VPWR VGND sg13g2_fill_1
X_2760_ _1005_ VPWR _1006_ VGND net836 _0601_ sg13g2_o21ai_1
XFILLER_8_552 VPWR VGND sg13g2_fill_1
X_2691_ net931 net556 _0954_ VPWR VGND sg13g2_nor2_1
X_4430_ net699 VGND VPWR _0421_ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
X_4361_ net641 VGND VPWR net912 net26 clknet_leaf_11_clk sg13g2_dfrbpq_2
X_4292_ net667 VGND VPWR net891 u_usb_cdc.u_ctrl_endp.max_length_q\[6\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
X_3312_ _1367_ net795 _1358_ VPWR VGND sg13g2_nand2_1
X_3243_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[19\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[27\]
+ net812 _1312_ VPWR VGND sg13g2_mux2_1
XFILLER_39_401 VPWR VGND sg13g2_decap_4
XFILLER_6_1024 VPWR VGND sg13g2_decap_4
X_3174_ _1248_ _1249_ _1250_ VPWR VGND sg13g2_nor2_1
X_2125_ net312 net210 _0060_ _2003_ VPWR VGND sg13g2_nand3_1
XFILLER_26_117 VPWR VGND sg13g2_fill_2
X_2056_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\] _1935_ VPWR VGND sg13g2_inv_4
XFILLER_35_695 VPWR VGND sg13g2_fill_1
XFILLER_10_518 VPWR VGND sg13g2_decap_8
X_2958_ net448 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ _1121_ _0151_ VPWR VGND sg13g2_mux2_1
X_2889_ _1096_ VPWR _0106_ VGND net824 _1097_ sg13g2_o21ai_1
Xhold530 _0027_ VPWR VGND net848 sg13g2_dlygate4sd3_1
Xhold552 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[1\] VPWR VGND
+ net870 sg13g2_dlygate4sd3_1
XFILLER_2_739 VPWR VGND sg13g2_decap_8
Xhold541 _0359_ VPWR VGND net859 sg13g2_dlygate4sd3_1
Xhold563 u_usb_cdc.u_sie.crc16_q\[8\] VPWR VGND net881 sg13g2_dlygate4sd3_1
Xhold585 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\] VPWR VGND
+ net903 sg13g2_dlygate4sd3_1
Xhold596 _0408_ VPWR VGND net914 sg13g2_dlygate4sd3_1
Xhold574 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[1\] VPWR VGND net892 sg13g2_dlygate4sd3_1
XFILLER_46_949 VPWR VGND sg13g2_decap_8
XFILLER_45_426 VPWR VGND sg13g2_fill_2
XFILLER_26_651 VPWR VGND sg13g2_fill_1
XFILLER_41_643 VPWR VGND sg13g2_fill_2
XFILLER_25_161 VPWR VGND sg13g2_fill_2
XFILLER_22_890 VPWR VGND sg13g2_decap_4
XFILLER_12_1007 VPWR VGND sg13g2_decap_8
XFILLER_31_83 VPWR VGND sg13g2_decap_4
XFILLER_1_750 VPWR VGND sg13g2_decap_8
XFILLER_49_732 VPWR VGND sg13g2_decap_8
XFILLER_45_982 VPWR VGND sg13g2_decap_8
X_3930_ _1823_ _1822_ _1817_ _1818_ net211 VPWR VGND sg13g2_a22oi_1
X_3861_ _1778_ VPWR _0395_ VGND _1779_ _1780_ sg13g2_o21ai_1
X_2812_ _1052_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[3\] _1053_
+ VPWR VGND sg13g2_xor2_1
X_3792_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] _0056_ _1728_ VPWR VGND sg13g2_nor2b_1
X_2743_ u_usb_cdc.u_ctrl_endp.state_q\[2\] u_usb_cdc.u_ctrl_endp.state_q\[6\] _0557_
+ _0748_ _0990_ VPWR VGND sg13g2_nor4_1
X_2674_ _0942_ net515 _0443_ VPWR VGND sg13g2_nand2_1
X_4413_ net729 VGND VPWR _0412_ u_usb_cdc.u_sie.rx_data\[0\] clknet_leaf_33_clk sg13g2_dfrbpq_2
X_4344_ net686 VGND VPWR _0346_ u_usb_cdc.u_sie.data_q\[7\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4275_ net693 VGND VPWR _0277_ u_usb_cdc.u_ctrl_endp.addr_dd\[2\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_3226_ _1297_ _1296_ net145 net601 net894 VPWR VGND sg13g2_a22oi_1
X_3157_ _1236_ net134 _1230_ VPWR VGND sg13g2_nand2_1
XFILLER_27_415 VPWR VGND sg13g2_decap_8
XFILLER_43_908 VPWR VGND sg13g2_decap_8
X_2108_ u_usb_cdc.endp\[1\] u_usb_cdc.endp\[3\] u_usb_cdc.endp\[2\] _1986_ VPWR VGND
+ sg13g2_nor3_2
XFILLER_42_407 VPWR VGND sg13g2_fill_1
X_3088_ _1199_ net98 _1193_ VPWR VGND sg13g2_nand2_1
XFILLER_36_982 VPWR VGND sg13g2_decap_8
X_2039_ VPWR _1918_ u_usb_cdc.u_ctrl_endp.req_q\[2\] VGND sg13g2_inv_1
XFILLER_10_326 VPWR VGND sg13g2_fill_1
XFILLER_2_536 VPWR VGND sg13g2_decap_8
Xhold360 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[8\] VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold371 u_usb_cdc.u_sie.phy_state_q\[2\] VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold382 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[2\] VPWR VGND
+ net424 sg13g2_dlygate4sd3_1
Xhold393 _0140_ VPWR VGND net435 sg13g2_dlygate4sd3_1
Xfanout840 net1050 net840 VPWR VGND sg13g2_buf_1
XFILLER_46_746 VPWR VGND sg13g2_decap_8
XFILLER_18_448 VPWR VGND sg13g2_fill_1
XFILLER_18_459 VPWR VGND sg13g2_decap_8
XFILLER_33_407 VPWR VGND sg13g2_decap_4
XFILLER_14_632 VPWR VGND sg13g2_fill_1
XFILLER_42_963 VPWR VGND sg13g2_decap_8
XFILLER_13_120 VPWR VGND sg13g2_fill_1
XFILLER_6_842 VPWR VGND sg13g2_decap_8
XFILLER_5_330 VPWR VGND sg13g2_fill_1
XFILLER_5_374 VPWR VGND sg13g2_decap_8
X_2390_ net587 net583 net619 _0689_ _0690_ VPWR VGND sg13g2_nor4_1
XFILLER_49_540 VPWR VGND sg13g2_decap_8
X_4060_ net728 VGND VPWR net258 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[4\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_49_584 VPWR VGND sg13g2_decap_8
X_3011_ net823 _1150_ net761 _1151_ VPWR VGND sg13g2_nand3_1
XFILLER_37_724 VPWR VGND sg13g2_decap_8
XFILLER_37_768 VPWR VGND sg13g2_decap_8
XFILLER_36_245 VPWR VGND sg13g2_decap_4
XFILLER_36_256 VPWR VGND sg13g2_fill_1
XFILLER_45_790 VPWR VGND sg13g2_decap_8
XFILLER_17_470 VPWR VGND sg13g2_decap_4
XFILLER_17_492 VPWR VGND sg13g2_decap_8
X_3913_ _1807_ _1805_ _1806_ VPWR VGND sg13g2_nand2_1
X_3844_ net303 _1765_ _1768_ VPWR VGND sg13g2_and2_1
XFILLER_20_624 VPWR VGND sg13g2_fill_2
XFILLER_20_657 VPWR VGND sg13g2_fill_1
X_3775_ _1718_ _0938_ _1936_ _0443_ net515 VPWR VGND sg13g2_a22oi_1
X_2726_ net48 net51 _0040_ VPWR VGND sg13g2_xor2_1
X_2657_ _0926_ VPWR _0927_ VGND _0700_ _0769_ sg13g2_o21ai_1
X_2588_ net745 _0498_ _0870_ VPWR VGND sg13g2_nor2_1
X_4327_ net688 VGND VPWR _0329_ u_usb_cdc.u_sie.crc16_q\[6\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_4258_ net683 VGND VPWR net1028 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[1\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3209_ net815 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[16\]
+ _1281_ VPWR VGND sg13g2_nor2_1
X_4189_ net665 VGND VPWR _0192_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[25\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_15_407 VPWR VGND sg13g2_decap_8
XFILLER_42_237 VPWR VGND sg13g2_fill_2
XFILLER_24_996 VPWR VGND sg13g2_decap_8
XFILLER_12_63 VPWR VGND sg13g2_fill_2
XFILLER_3_801 VPWR VGND sg13g2_decap_8
XFILLER_3_878 VPWR VGND sg13g2_decap_8
XFILLER_2_399 VPWR VGND sg13g2_decap_8
Xhold190 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[5\] VPWR VGND
+ net232 sg13g2_dlygate4sd3_1
Xfanout681 net682 net681 VPWR VGND sg13g2_buf_8
Xfanout692 net700 net692 VPWR VGND sg13g2_buf_2
Xfanout670 net671 net670 VPWR VGND sg13g2_buf_8
XFILLER_19_757 VPWR VGND sg13g2_fill_2
XFILLER_41_281 VPWR VGND sg13g2_fill_1
XFILLER_30_977 VPWR VGND sg13g2_decap_8
X_3560_ _1534_ VPWR _1535_ VGND net797 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[33\]
+ sg13g2_o21ai_1
X_2511_ net884 _0734_ _0736_ _0807_ _0808_ VPWR VGND sg13g2_nor4_1
X_3491_ _1482_ _0905_ _0595_ _1483_ VPWR VGND sg13g2_a21o_1
X_2442_ net860 _0739_ _0740_ VPWR VGND sg13g2_nor2_1
X_2373_ _0673_ _0672_ VPWR VGND _0649_ sg13g2_nand2b_2
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
X_4112_ net654 VGND VPWR net437 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[32\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4043_ net685 VGND VPWR net889 u_usb_cdc.u_ctrl_endp.state_q\[7\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_2
XFILLER_37_510 VPWR VGND sg13g2_fill_2
XFILLER_25_727 VPWR VGND sg13g2_decap_8
XFILLER_24_237 VPWR VGND sg13g2_decap_4
XFILLER_33_18 VPWR VGND sg13g2_decap_4
X_3827_ net278 _1747_ net740 _1756_ VPWR VGND sg13g2_nand3_1
XFILLER_20_487 VPWR VGND sg13g2_fill_1
X_3758_ _1704_ net833 _1703_ VPWR VGND sg13g2_nand2b_1
X_2709_ _0967_ net533 net11 VPWR VGND sg13g2_nand2b_1
X_3689_ _1646_ VPWR _1659_ VGND u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\]
+ _1658_ sg13g2_o21ai_1
XFILLER_0_815 VPWR VGND sg13g2_decap_8
XFILLER_48_819 VPWR VGND sg13g2_decap_8
XFILLER_28_543 VPWR VGND sg13g2_decap_8
XFILLER_12_944 VPWR VGND sg13g2_decap_8
XFILLER_11_443 VPWR VGND sg13g2_fill_1
XFILLER_23_62 VPWR VGND sg13g2_decap_4
XFILLER_8_959 VPWR VGND sg13g2_decap_8
XFILLER_11_476 VPWR VGND sg13g2_decap_4
XFILLER_3_675 VPWR VGND sg13g2_decap_8
XFILLER_39_808 VPWR VGND sg13g2_fill_2
XFILLER_47_863 VPWR VGND sg13g2_decap_8
XFILLER_19_565 VPWR VGND sg13g2_fill_1
XFILLER_19_576 VPWR VGND sg13g2_decap_8
X_2991_ _1138_ VPWR _0167_ VGND net721 _1137_ sg13g2_o21ai_1
XFILLER_14_281 VPWR VGND sg13g2_decap_8
XFILLER_9_75 VPWR VGND sg13g2_fill_2
XFILLER_30_763 VPWR VGND sg13g2_decap_4
X_3612_ VGND VPWR net800 _1970_ _1585_ net791 sg13g2_a21oi_1
XFILLER_30_796 VPWR VGND sg13g2_decap_4
XFILLER_31_1010 VPWR VGND sg13g2_decap_8
X_3543_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[1\] net779 _0547_ _1519_ VPWR VGND sg13g2_nor3_2
XFILLER_43_0 VPWR VGND sg13g2_fill_2
X_3474_ net460 _1471_ _1472_ VPWR VGND sg13g2_nor2_1
XFILLER_9_1022 VPWR VGND sg13g2_decap_8
X_2425_ net588 net585 _0682_ _0723_ VPWR VGND sg13g2_nor3_1
X_2356_ _0656_ _0655_ VPWR VGND sg13g2_inv_2
X_2287_ net746 net748 u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq _0589_ VPWR VGND sg13g2_nor3_2
XFILLER_38_830 VPWR VGND sg13g2_fill_1
X_4026_ net676 VGND VPWR net907 u_usb_cdc.u_ctrl_endp.req_q\[6\] clknet_leaf_47_clk
+ sg13g2_dfrbpq_2
XFILLER_44_28 VPWR VGND sg13g2_fill_2
XFILLER_13_708 VPWR VGND sg13g2_decap_8
XFILLER_25_557 VPWR VGND sg13g2_decap_8
XFILLER_20_262 VPWR VGND sg13g2_decap_4
XFILLER_5_918 VPWR VGND sg13g2_decap_8
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_0_612 VPWR VGND sg13g2_decap_8
XFILLER_48_627 VPWR VGND sg13g2_fill_1
XFILLER_0_689 VPWR VGND sg13g2_decap_8
XFILLER_28_351 VPWR VGND sg13g2_decap_8
XFILLER_44_822 VPWR VGND sg13g2_decap_8
XFILLER_44_899 VPWR VGND sg13g2_decap_8
XFILLER_31_538 VPWR VGND sg13g2_decap_8
XFILLER_15_1005 VPWR VGND sg13g2_decap_8
XFILLER_34_94 VPWR VGND sg13g2_fill_2
XFILLER_4_984 VPWR VGND sg13g2_decap_8
X_2210_ _0512_ _0510_ _0511_ VPWR VGND sg13g2_xnor2_1
X_3190_ _1264_ net768 net983 VPWR VGND sg13g2_nand2_1
XFILLER_15_4 VPWR VGND sg13g2_decap_4
X_2141_ VPWR _0444_ _0443_ VGND sg13g2_inv_1
X_2072_ _1951_ net285 VPWR VGND sg13g2_inv_2
XFILLER_34_376 VPWR VGND sg13g2_decap_4
X_2974_ _1049_ net825 _1055_ _0161_ VPWR VGND sg13g2_mux2_1
XFILLER_34_398 VPWR VGND sg13g2_fill_1
XFILLER_30_571 VPWR VGND sg13g2_decap_4
Xhold712 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[4\] VPWR VGND net1030 sg13g2_dlygate4sd3_1
Xhold701 _0369_ VPWR VGND net1019 sg13g2_dlygate4sd3_1
Xhold745 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[0\] VPWR VGND net1063 sg13g2_dlygate4sd3_1
X_3526_ net773 net770 _1502_ VPWR VGND sg13g2_nor2b_1
Xhold723 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ VPWR VGND net1041 sg13g2_dlygate4sd3_1
Xhold734 u_usb_cdc.u_sie.data_q\[1\] VPWR VGND net1052 sg13g2_dlygate4sd3_1
X_3457_ VGND VPWR _1457_ _1458_ _1459_ net878 sg13g2_a21oi_1
X_2408_ u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\]
+ u_usb_cdc.configured_o VPWR VGND sg13g2_and2_1
X_3388_ net756 _1408_ _1413_ VPWR VGND sg13g2_nor2_1
X_2339_ VGND VPWR u_usb_cdc.sie_in_req net634 _0640_ u_usb_cdc.sie_in_data_ack sg13g2_a21oi_1
XFILLER_45_619 VPWR VGND sg13g2_fill_1
X_4009_ _1887_ net634 _1884_ VPWR VGND sg13g2_nand2_1
XFILLER_38_1005 VPWR VGND sg13g2_decap_8
XFILLER_41_825 VPWR VGND sg13g2_decap_8
XFILLER_26_888 VPWR VGND sg13g2_fill_2
XFILLER_9_509 VPWR VGND sg13g2_decap_8
XFILLER_5_715 VPWR VGND sg13g2_decap_8
XFILLER_1_932 VPWR VGND sg13g2_decap_8
XFILLER_49_914 VPWR VGND sg13g2_decap_8
Xhold50 _0098_ VPWR VGND net92 sg13g2_dlygate4sd3_1
XFILLER_0_486 VPWR VGND sg13g2_decap_8
XFILLER_29_61 VPWR VGND sg13g2_fill_2
Xhold83 _0133_ VPWR VGND net125 sg13g2_dlygate4sd3_1
Xhold72 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[49\] VPWR VGND
+ net114 sg13g2_dlygate4sd3_1
Xhold61 _0178_ VPWR VGND net103 sg13g2_dlygate4sd3_1
Xhold94 _0052_ VPWR VGND net136 sg13g2_dlygate4sd3_1
XFILLER_29_671 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_55_clk clknet_3_0__leaf_clk clknet_leaf_55_clk VPWR VGND sg13g2_buf_8
XFILLER_17_855 VPWR VGND sg13g2_fill_2
XFILLER_44_652 VPWR VGND sg13g2_decap_8
XFILLER_16_376 VPWR VGND sg13g2_decap_4
XFILLER_43_195 VPWR VGND sg13g2_fill_1
XFILLER_8_531 VPWR VGND sg13g2_fill_2
X_2690_ net621 _2005_ _0953_ VPWR VGND sg13g2_nor2_1
X_4360_ net648 VGND VPWR net844 net21 clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3311_ _1365_ VPWR _1366_ VGND net927 _1128_ sg13g2_o21ai_1
XFILLER_4_781 VPWR VGND sg13g2_decap_8
XFILLER_3_280 VPWR VGND sg13g2_fill_1
X_4291_ net663 VGND VPWR net855 u_usb_cdc.u_ctrl_endp.max_length_q\[5\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_6_1003 VPWR VGND sg13g2_decap_8
X_3242_ VGND VPWR net809 _1306_ _1311_ _1310_ sg13g2_a21oi_1
X_3173_ _1249_ _1243_ _1148_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_435 VPWR VGND sg13g2_fill_2
X_2124_ _2002_ _0060_ net312 _0058_ VPWR VGND sg13g2_and3_2
XFILLER_48_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_46_clk clknet_3_5__leaf_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
X_2055_ _1934_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] VPWR VGND sg13g2_inv_2
X_2957_ net477 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ _1121_ _0150_ VPWR VGND sg13g2_mux2_1
X_2888_ _1097_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ _1082_ VPWR VGND sg13g2_nand2_1
Xhold520 _0958_ VPWR VGND net562 sg13g2_dlygate4sd3_1
Xhold542 _0048_ VPWR VGND net860 sg13g2_dlygate4sd3_1
XFILLER_2_718 VPWR VGND sg13g2_decap_8
Xhold553 u_usb_cdc.u_ctrl_endp.state_q\[3\] VPWR VGND net871 sg13g2_dlygate4sd3_1
Xhold531 u_usb_cdc.u_sie.out_toggle_q\[1\] VPWR VGND net849 sg13g2_dlygate4sd3_1
Xhold564 u_usb_cdc.u_sie.crc16_q\[7\] VPWR VGND net882 sg13g2_dlygate4sd3_1
Xhold597 u_usb_cdc.u_sie.crc16_q\[15\] VPWR VGND net915 sg13g2_dlygate4sd3_1
X_3509_ _1486_ _1952_ _1485_ VPWR VGND sg13g2_xnor2_1
Xhold575 _0029_ VPWR VGND net893 sg13g2_dlygate4sd3_1
Xhold586 u_usb_cdc.u_sie.pid_q\[0\] VPWR VGND net904 sg13g2_dlygate4sd3_1
XFILLER_46_928 VPWR VGND sg13g2_decap_8
XFILLER_39_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_37_clk clknet_3_5__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_26_663 VPWR VGND sg13g2_fill_1
XFILLER_41_622 VPWR VGND sg13g2_decap_8
XFILLER_13_335 VPWR VGND sg13g2_fill_2
Xoutput40 net40 usb_dp_tx_o VPWR VGND sg13g2_buf_1
XFILLER_49_711 VPWR VGND sg13g2_decap_8
XFILLER_49_788 VPWR VGND sg13g2_decap_8
XFILLER_48_276 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_28_clk clknet_3_7__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_36_438 VPWR VGND sg13g2_fill_2
XFILLER_45_961 VPWR VGND sg13g2_decap_8
XFILLER_44_493 VPWR VGND sg13g2_decap_8
X_3860_ _1739_ VPWR _1780_ VGND net297 _1776_ sg13g2_o21ai_1
X_2811_ _1044_ _1048_ _1052_ VPWR VGND sg13g2_and2_1
X_3791_ VPWR _0378_ net909 VGND sg13g2_inv_1
X_2742_ VPWR VGND _0988_ net170 _0985_ _1903_ _0067_ _0983_ sg13g2_a221oi_1
XFILLER_9_873 VPWR VGND sg13g2_decap_8
X_2673_ _0941_ VPWR _0030_ VGND _0934_ _0935_ sg13g2_o21ai_1
X_4412_ net729 VGND VPWR net530 u_usb_cdc.u_sie.u_phy_rx.rx_valid_q clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_28_1026 VPWR VGND sg13g2_fill_2
X_4343_ net686 VGND VPWR _0345_ u_usb_cdc.u_sie.data_q\[6\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4274_ net679 VGND VPWR _0276_ u_usb_cdc.u_ctrl_endp.addr_dd\[1\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
X_3225_ _1274_ _1287_ _1296_ VPWR VGND sg13g2_and2_1
X_3156_ _1235_ VPWR _0235_ VGND _1176_ _1229_ sg13g2_o21ai_1
Xclkbuf_leaf_19_clk clknet_3_3__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
X_3087_ _1198_ VPWR _0203_ VGND _1899_ net606 sg13g2_o21ai_1
X_2107_ VGND VPWR _1985_ u_usb_cdc.endp\[2\] u_usb_cdc.endp\[1\] sg13g2_or2_1
X_2038_ _1917_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] VPWR VGND sg13g2_inv_2
XFILLER_36_961 VPWR VGND sg13g2_decap_8
XFILLER_22_143 VPWR VGND sg13g2_fill_2
XFILLER_11_839 VPWR VGND sg13g2_fill_2
XFILLER_23_677 VPWR VGND sg13g2_fill_2
X_3989_ _1873_ _1033_ _1872_ net622 net1000 VPWR VGND sg13g2_a22oi_1
Xhold350 u_usb_cdc.u_ctrl_endp.addr_dd\[2\] VPWR VGND net392 sg13g2_dlygate4sd3_1
Xhold361 _0389_ VPWR VGND net403 sg13g2_dlygate4sd3_1
Xhold383 _0085_ VPWR VGND net425 sg13g2_dlygate4sd3_1
Xhold372 _0021_ VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold394 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[32\] VPWR VGND
+ net436 sg13g2_dlygate4sd3_1
Xfanout841 u_usb_cdc.u_ctrl_endp.state_q\[3\] net841 VPWR VGND sg13g2_buf_8
Xfanout830 u_usb_cdc.u_sie.phy_state_q\[11\] net830 VPWR VGND sg13g2_buf_8
XFILLER_46_725 VPWR VGND sg13g2_decap_8
XFILLER_19_917 VPWR VGND sg13g2_fill_2
XFILLER_27_983 VPWR VGND sg13g2_fill_2
XFILLER_42_942 VPWR VGND sg13g2_decap_8
XFILLER_13_187 VPWR VGND sg13g2_fill_2
XFILLER_6_821 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_fill_1
XFILLER_6_898 VPWR VGND sg13g2_decap_8
XFILLER_3_66 VPWR VGND sg13g2_fill_2
X_3010_ _1150_ net735 _1962_ _1149_ VPWR VGND sg13g2_and3_2
XFILLER_32_441 VPWR VGND sg13g2_decap_8
X_3912_ _1806_ _0585_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] _2003_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_3843_ _1767_ net710 net303 VPWR VGND sg13g2_nand2_1
XFILLER_32_463 VPWR VGND sg13g2_fill_2
XFILLER_33_986 VPWR VGND sg13g2_decap_8
X_3774_ VGND VPWR _1465_ _1710_ _0371_ net292 sg13g2_a21oi_1
X_2725_ VGND VPWR _0054_ net40 _1975_ net829 sg13g2_a21oi_2
X_2656_ _0693_ _0743_ _0675_ _0926_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_8_clk clknet_3_3__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_2587_ _0496_ net590 _0494_ _0869_ VPWR VGND _0601_ sg13g2_nand4_1
X_4326_ net687 VGND VPWR _0328_ u_usb_cdc.u_sie.crc16_q\[5\] clknet_leaf_27_clk sg13g2_dfrbpq_1
X_4257_ net683 VGND VPWR net1047 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[0\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_47_28 VPWR VGND sg13g2_fill_2
XFILLER_47_17 VPWR VGND sg13g2_decap_8
X_3208_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[0\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[8\]
+ net815 _1280_ VPWR VGND sg13g2_mux2_1
X_4188_ net665 VGND VPWR net228 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[24\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_3139_ _1226_ net167 net628 VPWR VGND sg13g2_nand2_1
XFILLER_28_736 VPWR VGND sg13g2_fill_2
XFILLER_42_216 VPWR VGND sg13g2_decap_4
XFILLER_27_279 VPWR VGND sg13g2_decap_4
XFILLER_24_942 VPWR VGND sg13g2_fill_1
XFILLER_24_975 VPWR VGND sg13g2_decap_8
XFILLER_3_857 VPWR VGND sg13g2_decap_8
Xhold180 _0182_ VPWR VGND net222 sg13g2_dlygate4sd3_1
XFILLER_2_378 VPWR VGND sg13g2_decap_8
Xhold191 _0172_ VPWR VGND net233 sg13g2_dlygate4sd3_1
Xfanout660 net661 net660 VPWR VGND sg13g2_buf_2
Xfanout693 net700 net693 VPWR VGND sg13g2_buf_8
Xfanout682 net690 net682 VPWR VGND sg13g2_buf_8
Xfanout671 net675 net671 VPWR VGND sg13g2_buf_8
XFILLER_18_257 VPWR VGND sg13g2_fill_1
XFILLER_19_769 VPWR VGND sg13g2_decap_4
XFILLER_15_920 VPWR VGND sg13g2_decap_8
XFILLER_18_1014 VPWR VGND sg13g2_decap_8
XFILLER_30_956 VPWR VGND sg13g2_decap_8
X_2510_ _0797_ _0804_ _0805_ _0806_ _0807_ VPWR VGND sg13g2_nor4_1
X_3490_ net834 net839 net836 _1482_ VPWR VGND sg13g2_nor3_1
X_2441_ _0653_ _0738_ net736 _0739_ VPWR VGND sg13g2_nand3_1
X_2372_ _0666_ _0668_ _0669_ _0671_ _0672_ VPWR VGND sg13g2_nor4_1
X_4111_ net668 VGND VPWR net474 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[31\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_4042_ net678 VGND VPWR net1004 u_usb_cdc.u_ctrl_endp.state_q\[6\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_2
XFILLER_49_382 VPWR VGND sg13g2_fill_2
XFILLER_20_422 VPWR VGND sg13g2_decap_4
X_3826_ net712 _1754_ _1755_ VPWR VGND sg13g2_nor2_1
X_3757_ _1703_ net633 net769 _0572_ u_usb_cdc.ctrl_stall VPWR VGND sg13g2_a22oi_1
X_2708_ net735 VPWR _0966_ VGND _0963_ _0965_ sg13g2_o21ai_1
X_3688_ _1651_ VPWR _1658_ VGND _1654_ _1657_ sg13g2_o21ai_1
X_2639_ VPWR _0019_ _0910_ VGND sg13g2_inv_1
X_4309_ net693 VGND VPWR net215 u_usb_cdc.u_sie.addr_q\[5\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_28_533 VPWR VGND sg13g2_fill_1
XFILLER_12_923 VPWR VGND sg13g2_decap_8
XFILLER_11_411 VPWR VGND sg13g2_decap_8
XFILLER_23_260 VPWR VGND sg13g2_decap_8
XFILLER_24_783 VPWR VGND sg13g2_fill_1
XFILLER_8_938 VPWR VGND sg13g2_decap_8
XFILLER_23_41 VPWR VGND sg13g2_decap_8
XFILLER_11_499 VPWR VGND sg13g2_fill_1
XFILLER_3_654 VPWR VGND sg13g2_decap_8
XFILLER_47_842 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_fill_1
XFILLER_0_89 VPWR VGND sg13g2_fill_1
X_2990_ _1138_ net255 net613 VPWR VGND sg13g2_nand2_1
XFILLER_9_65 VPWR VGND sg13g2_fill_1
X_3611_ net797 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[3\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[11\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[19\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[27\]
+ net791 _1584_ VPWR VGND sg13g2_mux4_1
X_3542_ VGND VPWR _1514_ _1515_ _1518_ _1516_ sg13g2_a21oi_1
X_3473_ u_usb_cdc.u_sie.delay_cnt_q\[0\] net742 net507 _1471_ VPWR VGND sg13g2_nand3_1
XFILLER_9_1001 VPWR VGND sg13g2_decap_8
X_2424_ _0693_ _0713_ _0675_ _0722_ VPWR VGND sg13g2_nand3_1
X_2355_ _0655_ net784 _0653_ VPWR VGND sg13g2_nand2_2
X_2286_ _0585_ _0587_ _0588_ VPWR VGND sg13g2_nor2_1
X_4025_ net677 VGND VPWR _0006_ u_usb_cdc.u_ctrl_endp.req_q\[5\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
XFILLER_38_842 VPWR VGND sg13g2_fill_1
XFILLER_25_536 VPWR VGND sg13g2_decap_8
XFILLER_12_219 VPWR VGND sg13g2_fill_1
XFILLER_40_539 VPWR VGND sg13g2_decap_8
XFILLER_20_241 VPWR VGND sg13g2_fill_2
XFILLER_21_764 VPWR VGND sg13g2_fill_1
X_3809_ VGND VPWR net318 net331 _1742_ _1738_ sg13g2_a21oi_1
XFILLER_20_252 VPWR VGND sg13g2_decap_4
XFILLER_0_668 VPWR VGND sg13g2_decap_8
XFILLER_29_875 VPWR VGND sg13g2_fill_2
XFILLER_44_878 VPWR VGND sg13g2_decap_8
XFILLER_43_366 VPWR VGND sg13g2_fill_1
XFILLER_31_528 VPWR VGND sg13g2_decap_4
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_724 VPWR VGND sg13g2_decap_8
XFILLER_7_234 VPWR VGND sg13g2_fill_2
XFILLER_7_267 VPWR VGND sg13g2_decap_8
XFILLER_4_963 VPWR VGND sg13g2_decap_8
XFILLER_39_606 VPWR VGND sg13g2_decap_8
X_2140_ _2012_ _0440_ _0442_ _0443_ VPWR VGND sg13g2_nor3_2
X_2071_ _1950_ net306 VPWR VGND sg13g2_inv_2
X_2973_ _1045_ net827 _1055_ _0160_ VPWR VGND sg13g2_mux2_1
XFILLER_22_539 VPWR VGND sg13g2_fill_2
Xhold702 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] VPWR VGND
+ net1020 sg13g2_dlygate4sd3_1
Xhold735 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[1\] VPWR VGND
+ net1053 sg13g2_dlygate4sd3_1
Xhold746 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[3\] VPWR
+ VGND net1064 sg13g2_dlygate4sd3_1
Xhold713 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[5\] VPWR VGND net1031 sg13g2_dlygate4sd3_1
X_3525_ net625 VPWR _1501_ VGND _0576_ _1500_ sg13g2_o21ai_1
Xhold724 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ VPWR VGND net1042 sg13g2_dlygate4sd3_1
X_3456_ u_usb_cdc.u_ctrl_endp.req_q\[5\] u_usb_cdc.u_ctrl_endp.addr_dd\[1\] u_usb_cdc.u_ctrl_endp.addr_dd\[0\]
+ u_usb_cdc.u_ctrl_endp.addr_dd\[3\] _1458_ VPWR VGND sg13g2_nor4_1
X_2407_ _0061_ net574 _0706_ _0692_ _1982_ VPWR VGND sg13g2_a22oi_1
X_3387_ net523 net567 _1412_ VPWR VGND sg13g2_nor2_1
X_2338_ VGND VPWR _0639_ net583 net588 sg13g2_or2_1
X_2269_ _0563_ _0570_ _0571_ VPWR VGND sg13g2_nor2_1
X_4008_ _1886_ VPWR _0436_ VGND _1910_ _1885_ sg13g2_o21ai_1
XFILLER_25_344 VPWR VGND sg13g2_decap_4
XFILLER_26_878 VPWR VGND sg13g2_decap_4
XFILLER_40_369 VPWR VGND sg13g2_decap_8
XFILLER_1_911 VPWR VGND sg13g2_decap_8
XFILLER_1_988 VPWR VGND sg13g2_decap_8
Xhold40 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[2\] VPWR VGND
+ net82 sg13g2_dlygate4sd3_1
XFILLER_0_465 VPWR VGND sg13g2_decap_8
Xhold51 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[21\] VPWR VGND
+ net93 sg13g2_dlygate4sd3_1
Xhold62 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[8\] VPWR VGND
+ net104 sg13g2_dlygate4sd3_1
XFILLER_29_95 VPWR VGND sg13g2_fill_2
Xhold73 _0132_ VPWR VGND net115 sg13g2_dlygate4sd3_1
Xhold95 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[11\] VPWR VGND
+ net137 sg13g2_dlygate4sd3_1
Xhold84 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[52\] VPWR VGND
+ net126 sg13g2_dlygate4sd3_1
XFILLER_17_845 VPWR VGND sg13g2_fill_1
XFILLER_17_878 VPWR VGND sg13g2_fill_1
XFILLER_31_303 VPWR VGND sg13g2_fill_2
XFILLER_31_369 VPWR VGND sg13g2_decap_4
XFILLER_6_77 VPWR VGND sg13g2_decap_4
XFILLER_4_760 VPWR VGND sg13g2_decap_8
X_3310_ _1365_ _1128_ _1364_ VPWR VGND sg13g2_nand2_1
X_4290_ net663 VGND VPWR net539 u_usb_cdc.u_ctrl_endp.max_length_q\[4\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_3241_ net807 VPWR _1310_ VGND net809 _1308_ sg13g2_o21ai_1
X_3172_ VGND VPWR net820 _1183_ _1248_ net1017 sg13g2_a21oi_1
X_2123_ _2001_ net312 net210 VPWR VGND sg13g2_nand2_1
XFILLER_26_119 VPWR VGND sg13g2_fill_1
XFILLER_47_480 VPWR VGND sg13g2_decap_8
X_2054_ VPWR _1933_ net949 VGND sg13g2_inv_1
XFILLER_35_631 VPWR VGND sg13g2_decap_4
XFILLER_35_686 VPWR VGND sg13g2_decap_8
X_2956_ net464 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ _1121_ _0149_ VPWR VGND sg13g2_mux2_1
X_2887_ _1096_ net67 _1080_ VPWR VGND sg13g2_nand2_1
Xhold510 u_usb_cdc.u_ctrl_endp.req_q\[11\] VPWR VGND net552 sg13g2_dlygate4sd3_1
Xhold521 u_usb_cdc.u_sie.crc16_q\[13\] VPWR VGND net563 sg13g2_dlygate4sd3_1
Xhold543 _0061_ VPWR VGND net861 sg13g2_dlygate4sd3_1
Xhold554 _0013_ VPWR VGND net872 sg13g2_dlygate4sd3_1
Xhold532 _1002_ VPWR VGND net850 sg13g2_dlygate4sd3_1
Xhold565 _0330_ VPWR VGND net883 sg13g2_dlygate4sd3_1
X_3508_ _0337_ net573 _1953_ net576 _1939_ VPWR VGND sg13g2_a22oi_1
Xhold587 u_usb_cdc.addr\[3\] VPWR VGND net905 sg13g2_dlygate4sd3_1
Xhold576 net30 VPWR VGND net894 sg13g2_dlygate4sd3_1
Xhold598 u_usb_cdc.u_ctrl_endp.max_length_q\[3\] VPWR VGND net916 sg13g2_dlygate4sd3_1
X_3439_ net762 net582 _1448_ VPWR VGND sg13g2_nor2_1
XFILLER_46_907 VPWR VGND sg13g2_decap_8
XFILLER_18_609 VPWR VGND sg13g2_decap_8
XFILLER_25_163 VPWR VGND sg13g2_fill_1
XFILLER_41_667 VPWR VGND sg13g2_decap_4
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_13_358 VPWR VGND sg13g2_fill_1
XFILLER_15_53 VPWR VGND sg13g2_fill_1
XFILLER_25_196 VPWR VGND sg13g2_decap_4
XFILLER_15_86 VPWR VGND sg13g2_fill_2
Xoutput30 net30 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_785 VPWR VGND sg13g2_decap_8
XFILLER_49_767 VPWR VGND sg13g2_decap_8
XFILLER_45_940 VPWR VGND sg13g2_decap_8
X_2810_ _1044_ _1046_ _1042_ _1051_ VPWR VGND _1050_ sg13g2_nand4_1
X_3790_ _1727_ _1720_ net908 _0933_ net862 VPWR VGND sg13g2_a22oi_1
X_2741_ VGND VPWR _1906_ _0988_ _0989_ net169 sg13g2_a21oi_1
XFILLER_9_885 VPWR VGND sg13g2_decap_8
X_2672_ VPWR VGND net635 _0940_ _0938_ net1012 _0941_ net579 sg13g2_a221oi_1
X_4411_ net685 VGND VPWR net1035 u_usb_cdc.sie_in_data_ack clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_28_1005 VPWR VGND sg13g2_decap_8
X_4342_ net686 VGND VPWR _0344_ u_usb_cdc.u_sie.data_q\[5\] clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4273_ net679 VGND VPWR _0275_ u_usb_cdc.u_ctrl_endp.addr_dd\[0\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
X_3224_ net805 net601 _1294_ _1295_ VPWR VGND sg13g2_nor3_1
.ends

