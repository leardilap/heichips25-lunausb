VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spad_env_f_bit
  CLASS BLOCK ;
  FOREIGN spad_env_f_bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 21.580 3.560 23.780 68.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.660 22.480 72.220 24.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 15.380 3.560 17.580 68.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.660 16.280 72.220 18.480 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 18.700 0.400 19.100 ;
    END
  END clk
  PIN env_bit
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 74.600 18.700 75.000 19.100 ;
    END
  END env_bit
  PIN env_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 74.600 55.660 75.000 56.060 ;
    END
  END env_valid
  PIN spad_hit_async
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 55.660 0.400 56.060 ;
    END
  END spad_hit_async
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 72.000 68.190 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 72.000 68.260 ;
      LAYER Metal2 ;
        RECT 3.260 3.635 71.625 68.185 ;
      LAYER Metal3 ;
        RECT 0.400 56.270 74.600 68.140 ;
        RECT 0.610 55.450 74.390 56.270 ;
        RECT 0.400 19.310 74.600 55.450 ;
        RECT 0.610 18.490 74.390 19.310 ;
        RECT 0.400 3.680 74.600 18.490 ;
  END
END spad_env_f_bit
END LIBRARY

