module spad_env_f_bit (clk,
    env_bit,
    env_valid,
    spad_hit_async,
    VPWR,
    VGND);
 input clk;
 output env_bit;
 output env_valid;
 input spad_hit_async;
 inout VPWR;
 inout VGND;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire clknet_0_clk;
 wire net2;
 wire net3;
 wire prev2_bit;
 wire \pulse_cnt[0] ;
 wire \pulse_cnt[1] ;
 wire \pulse_cnt[2] ;
 wire \pulse_cnt[3] ;
 wire rise_spad;
 wire s0;
 wire s1;
 wire s1_d;
 wire \win_cnt[0] ;
 wire \win_cnt[10] ;
 wire \win_cnt[11] ;
 wire \win_cnt[12] ;
 wire \win_cnt[13] ;
 wire \win_cnt[14] ;
 wire \win_cnt[15] ;
 wire \win_cnt[1] ;
 wire \win_cnt[2] ;
 wire \win_cnt[3] ;
 wire \win_cnt[4] ;
 wire \win_cnt[5] ;
 wire \win_cnt[6] ;
 wire \win_cnt[7] ;
 wire \win_cnt[8] ;
 wire \win_cnt[9] ;
 wire win_rollover;
 wire net1;
 wire net4;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;

 sg13g2_inv_1 _082_ (.VDD(VPWR),
    .Y(_007_),
    .A(net36),
    .VSS(VGND));
 sg13g2_inv_1 _083_ (.VDD(VPWR),
    .Y(_025_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _084_ (.VDD(VPWR),
    .Y(_026_),
    .A(net41),
    .VSS(VGND));
 sg13g2_nand3_1 _085_ (.B(net72),
    .C(net76),
    .A(net36),
    .Y(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _086_ (.A(net36),
    .B(\win_cnt[1] ),
    .C(net39),
    .D(\win_cnt[2] ),
    .X(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _087_ (.A(net55),
    .B(_028_),
    .X(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _088_ (.B(net55),
    .C(net75),
    .A(net61),
    .Y(_030_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_028_));
 sg13g2_nor2_1 _089_ (.A(_025_),
    .B(_030_),
    .Y(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _090_ (.Y(_032_),
    .A(net48),
    .B(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _091_ (.A(_025_),
    .B(_030_),
    .C(_032_),
    .Y(_033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _092_ (.Y(_034_),
    .A(net43),
    .B(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _093_ (.A(_025_),
    .B(_030_),
    .C(_032_),
    .Y(_035_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_034_));
 sg13g2_nand3_1 _094_ (.B(net57),
    .C(_035_),
    .A(net51),
    .Y(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _095_ (.B(\win_cnt[12] ),
    .C(\win_cnt[14] ),
    .A(net51),
    .Y(_037_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_035_));
 sg13g2_nor2_1 _096_ (.A(_026_),
    .B(net52),
    .Y(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _097_ (.A(net34),
    .B_N(net33),
    .Y(_000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _098_ (.B(\pulse_cnt[2] ),
    .A(\pulse_cnt[3] ),
    .X(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _099_ (.Y(_039_),
    .A(\pulse_cnt[1] ),
    .B(\pulse_cnt[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _100_ (.Y(_040_),
    .A(_038_),
    .B(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _101_ (.B1(net35),
    .VDD(VPWR),
    .Y(_041_),
    .VSS(VGND),
    .A1(prev2_bit),
    .A2(_040_));
 sg13g2_a21oi_1 _102_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(prev2_bit),
    .A2(_040_),
    .Y(_042_),
    .B1(_041_));
 sg13g2_xor2_1 _103_ (.B(_042_),
    .A(net46),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _104_ (.Y(_043_),
    .A(rise_spad),
    .B(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _105_ (.A(net35),
    .B(net64),
    .Y(_003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _106_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(rise_spad),
    .A2(net63),
    .Y(_044_),
    .B1(net69));
 sg13g2_and3_1 _107_ (.X(_045_),
    .A(rise_spad),
    .B(net69),
    .C(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _108_ (.A(net35),
    .B(net70),
    .C(_045_),
    .Y(_004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _109_ (.A(net67),
    .B(_045_),
    .Y(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _110_ (.A(net67),
    .B(_045_),
    .X(_047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _111_ (.A(net35),
    .B(net68),
    .C(_047_),
    .Y(_005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _112_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net74),
    .A2(_047_),
    .Y(_048_),
    .B1(net35));
 sg13g2_o21ai_1 _113_ (.B1(_048_),
    .VDD(VPWR),
    .Y(_049_),
    .VSS(VGND),
    .A1(net74),
    .A2(_047_));
 sg13g2_inv_1 _114_ (.VDD(VPWR),
    .Y(_006_),
    .A(_049_),
    .VSS(VGND));
 sg13g2_xor2_1 _115_ (.B(net72),
    .A(net36),
    .X(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _116_ (.A2(net72),
    .A1(net36),
    .B1(net76),
    .X(_050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _117_ (.A(_027_),
    .B(_050_),
    .X(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _118_ (.Y(_010_),
    .A(net39),
    .B(_027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _119_ (.B(_028_),
    .A(net55),
    .X(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _120_ (.B(_029_),
    .A(net61),
    .X(_012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _121_ (.A2(_029_),
    .A1(net61),
    .B1(net75),
    .X(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _122_ (.A(_030_),
    .B(_051_),
    .X(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _123_ (.Y(_014_),
    .A(net37),
    .B(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _124_ (.B(_031_),
    .A(net59),
    .X(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _125_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\win_cnt[8] ),
    .A2(_031_),
    .Y(_052_),
    .B1(net48));
 sg13g2_nor2_1 _126_ (.A(_033_),
    .B(net49),
    .Y(_016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _127_ (.B(_033_),
    .A(net65),
    .X(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _128_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\win_cnt[10] ),
    .A2(_033_),
    .Y(_053_),
    .B1(net43));
 sg13g2_nor2_1 _129_ (.A(_035_),
    .B(net44),
    .Y(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _130_ (.B(_035_),
    .A(net57),
    .X(_019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _131_ (.A2(_035_),
    .A1(net57),
    .B1(net51),
    .X(_024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _132_ (.A(_036_),
    .B(_024_),
    .X(_020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _133_ (.Y(_021_),
    .A(net53),
    .B(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _134_ (.Y(_022_),
    .A(net41),
    .B(_037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _135_ (.A0(net73),
    .A1(net46),
    .S(net35),
    .X(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_2 _136_ (.RESET_B(net6),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net47),
    .Q(net2),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _137_ (.RESET_B(net7),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1),
    .Q(s0),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _138_ (.RESET_B(net8),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net32),
    .Q(s1),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _139_ (.RESET_B(net9),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net33),
    .Q(s1_d),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _140_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_000_),
    .Q(rise_spad),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _141_ (.RESET_B(net5),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_001_),
    .Q(win_rollover),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _142_ (.RESET_B(net20),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_003_),
    .Q(\pulse_cnt[0] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _143_ (.RESET_B(net18),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net71),
    .Q(\pulse_cnt[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _144_ (.RESET_B(net16),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_005_),
    .Q(\pulse_cnt[2] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _145_ (.RESET_B(net14),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_006_),
    .Q(\pulse_cnt[3] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _146_ (.RESET_B(net12),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_007_),
    .Q(\win_cnt[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _147_ (.RESET_B(net11),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_008_),
    .Q(\win_cnt[1] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _148_ (.RESET_B(net10),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_009_),
    .Q(\win_cnt[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _149_ (.RESET_B(net4),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net40),
    .Q(\win_cnt[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _150_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net56),
    .Q(\win_cnt[4] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _151_ (.RESET_B(net29),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net62),
    .Q(\win_cnt[5] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _152_ (.RESET_B(net28),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_013_),
    .Q(\win_cnt[6] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _153_ (.RESET_B(net27),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net38),
    .Q(\win_cnt[7] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _154_ (.RESET_B(net26),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net60),
    .Q(\win_cnt[8] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _155_ (.RESET_B(net25),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net50),
    .Q(\win_cnt[9] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _156_ (.RESET_B(net24),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net66),
    .Q(\win_cnt[10] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _157_ (.RESET_B(net23),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net45),
    .Q(\win_cnt[11] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _158_ (.RESET_B(net22),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net58),
    .Q(\win_cnt[12] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _159_ (.RESET_B(net21),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_020_),
    .Q(\win_cnt[13] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _160_ (.RESET_B(net19),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net54),
    .Q(\win_cnt[14] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _161_ (.RESET_B(net17),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net42),
    .Q(\win_cnt[15] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _162_ (.RESET_B(net13),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_023_),
    .Q(prev2_bit),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _163_ (.RESET_B(net15),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net35),
    .Q(net3),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_tiehi _141__5 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net5));
 sg13g2_tiehi _136__6 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net6));
 sg13g2_tiehi _137__7 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net7));
 sg13g2_tiehi _138__8 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net8));
 sg13g2_tiehi _139__9 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net9));
 sg13g2_tiehi _148__10 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net10));
 sg13g2_tiehi _147__11 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net11));
 sg13g2_tiehi _146__12 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net12));
 sg13g2_tiehi _162__13 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net13));
 sg13g2_tiehi _145__14 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net14));
 sg13g2_tiehi _163__15 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net15));
 sg13g2_tiehi _144__16 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net16));
 sg13g2_tiehi _161__17 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net17));
 sg13g2_tiehi _143__18 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net18));
 sg13g2_tiehi _160__19 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net19));
 sg13g2_tiehi _142__20 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net20));
 sg13g2_tiehi _159__21 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net21));
 sg13g2_tiehi _158__22 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net22));
 sg13g2_tiehi _157__23 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net23));
 sg13g2_tiehi _156__24 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net24));
 sg13g2_tiehi _155__25 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net25));
 sg13g2_tiehi _154__26 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net26));
 sg13g2_tiehi _153__27 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net27));
 sg13g2_tiehi _152__28 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net28));
 sg13g2_tiehi _151__29 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net29));
 sg13g2_tiehi _150__30 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net30));
 sg13g2_tiehi _140__31 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net31));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(spad_hit_async),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(env_bit),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(env_valid),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _149__4 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net4));
 sg13g2_buf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload0 (.A(clknet_2_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload1 (.A(clknet_2_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(s0),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold2 (.A(s1),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold3 (.A(s1_d),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold4 (.A(win_rollover),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold5 (.A(\win_cnt[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold6 (.A(\win_cnt[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold7 (.A(_014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold8 (.A(\win_cnt[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold9 (.A(_010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold10 (.A(\win_cnt[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold11 (.A(_022_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold12 (.A(\win_cnt[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold13 (.A(_053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold14 (.A(_018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold15 (.A(net2),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold16 (.A(_002_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold17 (.A(\win_cnt[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold18 (.A(_052_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold19 (.A(_016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold20 (.A(\win_cnt[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold21 (.A(_037_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold22 (.A(\win_cnt[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold23 (.A(_021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold24 (.A(\win_cnt[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold25 (.A(_011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold26 (.A(\win_cnt[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold27 (.A(_019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold28 (.A(\win_cnt[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold29 (.A(_015_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold30 (.A(\win_cnt[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold31 (.A(_012_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold32 (.A(\pulse_cnt[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold33 (.A(_043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold34 (.A(\win_cnt[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold35 (.A(_017_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold36 (.A(\pulse_cnt[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold37 (.A(_046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold38 (.A(\pulse_cnt[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold39 (.A(_044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold40 (.A(_004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold41 (.A(\win_cnt[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold42 (.A(prev2_bit),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold43 (.A(\pulse_cnt[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold44 (.A(\win_cnt[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold45 (.A(\win_cnt[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net76));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_142 (.VDD(VPWR),
    .VSS(VGND));
endmodule
