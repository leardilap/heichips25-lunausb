* NGSPICE file created from heichips25_usb_cdc.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for spad_env_f_bit abstract view
.subckt spad_env_f_bit VGND VPWR clk env_bit env_valid spad_hit_async
.ends

.subckt heichips25_usb_cdc VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] usb_dn_en_o usb_dn_rx_i usb_dn_tx_o usb_dp_en_o usb_dp_rx_i
+ usb_dp_tx_o usb_dp_up_o
X_3155_ _1202_ VPWR _0197_ VGND _1917_ net607 sg13g2_o21ai_1
X_3086_ net826 _1154_ net739 _1156_ VPWR VGND sg13g2_nand3_1
X_2106_ VPWR _1963_ net932 VGND sg13g2_inv_1
X_3988_ net754 _0925_ _1823_ VPWR VGND sg13g2_nor2_2
XFILLER_23_678 VPWR VGND sg13g2_fill_1
XFILLER_10_328 VPWR VGND sg13g2_decap_4
X_2939_ _1015_ net621 _1077_ VPWR VGND sg13g2_nor2_2
XFILLER_2_516 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_fill_2
Xhold340 u_usb_cdc.u_sie.u_phy_tx.data_q\[3\] VPWR VGND net383 sg13g2_dlygate4sd3_1
Xhold362 _0424_ VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold351 _0919_ VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold384 _0221_ VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold373 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[50\] VPWR
+ VGND net416 sg13g2_dlygate4sd3_1
Xhold395 _0381_ VPWR VGND net438 sg13g2_dlygate4sd3_1
Xfanout820 net1041 net820 VPWR VGND sg13g2_buf_8
Xfanout842 net843 net842 VPWR VGND sg13g2_buf_8
Xfanout831 net832 net831 VPWR VGND sg13g2_buf_1
XFILLER_46_704 VPWR VGND sg13g2_decap_8
XFILLER_27_951 VPWR VGND sg13g2_fill_1
XFILLER_42_910 VPWR VGND sg13g2_decap_8
XFILLER_42_987 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk_regs clknet_0_clk_regs clknet_3_6__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_49_520 VPWR VGND sg13g2_decap_8
XFILLER_49_597 VPWR VGND sg13g2_decap_8
X_3911_ net615 VPWR _1776_ VGND net340 _1772_ sg13g2_o21ai_1
X_3842_ _1726_ VPWR _1727_ VGND _0578_ _0956_ sg13g2_o21ai_1
XFILLER_33_998 VPWR VGND sg13g2_decap_8
X_3773_ _0439_ VPWR _1673_ VGND net506 _1523_ sg13g2_o21ai_1
X_2724_ net394 VPWR _0033_ VGND _1977_ _0917_ sg13g2_o21ai_1
X_2655_ _0843_ VPWR _0021_ VGND _0845_ _0865_ sg13g2_o21ai_1
X_4325_ net652 VGND VPWR net952 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[3\]
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_2
X_2586_ _0807_ net974 _0808_ _0009_ VPWR VGND sg13g2_a21o_1
X_4256_ net654 VGND VPWR net326 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[18\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_3207_ net396 net631 _1230_ VPWR VGND sg13g2_nor2_1
X_4187_ net667 VGND VPWR net219 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[33\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
X_3138_ VGND VPWR net633 _1192_ _0190_ net334 sg13g2_a21oi_1
XFILLER_27_214 VPWR VGND sg13g2_fill_2
X_3069_ _1145_ net288 net634 VPWR VGND sg13g2_nand2_1
XFILLER_24_998 VPWR VGND sg13g2_decap_8
XFILLER_6_129 VPWR VGND sg13g2_fill_2
XFILLER_3_847 VPWR VGND sg13g2_decap_4
Xhold170 _0206_ VPWR VGND net213 sg13g2_dlygate4sd3_1
XFILLER_2_379 VPWR VGND sg13g2_decap_8
Xhold192 _0213_ VPWR VGND net235 sg13g2_dlygate4sd3_1
Xhold181 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[56\] VPWR
+ VGND net224 sg13g2_dlygate4sd3_1
Xfanout650 net651 net650 VPWR VGND sg13g2_buf_2
Xfanout683 net685 net683 VPWR VGND sg13g2_buf_8
Xfanout672 net674 net672 VPWR VGND sg13g2_buf_8
Xfanout661 net665 net661 VPWR VGND sg13g2_buf_8
Xfanout694 net706 net694 VPWR VGND sg13g2_buf_8
XFILLER_15_965 VPWR VGND sg13g2_fill_2
XFILLER_30_968 VPWR VGND sg13g2_decap_8
X_2440_ _0670_ _1925_ net787 VPWR VGND sg13g2_nand2_1
X_2371_ _0601_ _0602_ VPWR VGND sg13g2_inv_4
XFILLER_38_4 VPWR VGND sg13g2_decap_8
X_4110_ net693 VGND VPWR net542 _0049_ clknet_leaf_33_clk_regs sg13g2_dfrbpq_1
X_4041_ _1865_ VPWR _0415_ VGND _1869_ _1870_ sg13g2_o21ai_1
XFILLER_49_394 VPWR VGND sg13g2_decap_8
X_3825_ _0990_ _1704_ _1712_ VPWR VGND sg13g2_nor2b_2
X_3756_ _1627_ VPWR _1657_ VGND _1628_ _1656_ sg13g2_o21ai_1
X_2707_ net976 _2038_ net1007 _0906_ VPWR VGND sg13g2_nand3_1
X_3687_ VGND VPWR net799 _1589_ _1590_ net796 sg13g2_a21oi_1
X_2638_ u_usb_cdc.u_sie.addr_q\[6\] u_usb_cdc.addr\[6\] _0849_ VPWR VGND sg13g2_xor2_1
X_2569_ VPWR VGND net588 _0792_ _0793_ _0663_ _0794_ net622 sg13g2_a221oi_1
X_4308_ net648 VGND VPWR net167 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[70\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
XFILLER_0_839 VPWR VGND sg13g2_fill_1
X_4239_ net675 VGND VPWR _0168_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[1\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
XFILLER_47_309 VPWR VGND sg13g2_decap_8
XFILLER_28_523 VPWR VGND sg13g2_fill_1
XFILLER_28_512 VPWR VGND sg13g2_fill_2
XFILLER_16_707 VPWR VGND sg13g2_fill_2
XFILLER_11_478 VPWR VGND sg13g2_decap_4
XFILLER_11_467 VPWR VGND sg13g2_fill_2
XFILLER_47_810 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_47_887 VPWR VGND sg13g2_decap_8
XFILLER_15_751 VPWR VGND sg13g2_fill_2
XFILLER_15_784 VPWR VGND sg13g2_fill_2
XFILLER_42_581 VPWR VGND sg13g2_fill_1
X_3610_ _0545_ VPWR _1516_ VGND _1514_ _1515_ sg13g2_o21ai_1
XFILLER_31_1023 VPWR VGND sg13g2_decap_4
X_3541_ _1469_ VPWR _1472_ VGND _1940_ net179 sg13g2_o21ai_1
XFILLER_7_972 VPWR VGND sg13g2_decap_8
X_3472_ VGND VPWR net576 _1426_ _0290_ _1425_ sg13g2_a21oi_1
XFILLER_9_1002 VPWR VGND sg13g2_decap_8
X_2423_ _0540_ net785 net781 _0653_ VPWR VGND sg13g2_a21o_1
X_2354_ u_usb_cdc.u_sie.in_byte_q\[3\] _2017_ _0584_ _0585_ VPWR VGND sg13g2_nor3_1
X_2285_ _0517_ u_usb_cdc.ctrl_stall net640 VPWR VGND sg13g2_nand2_1
X_4024_ _2027_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] _1830_ _1856_ VPWR VGND sg13g2_a21o_1
X_3808_ _1699_ VPWR _0353_ VGND _1917_ net600 sg13g2_o21ai_1
X_3739_ VGND VPWR net804 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[13\]
+ _1640_ _1639_ sg13g2_a21oi_1
XFILLER_0_636 VPWR VGND sg13g2_decap_8
XFILLER_44_879 VPWR VGND sg13g2_decap_8
XFILLER_12_732 VPWR VGND sg13g2_fill_1
XFILLER_12_787 VPWR VGND sg13g2_fill_1
XFILLER_4_953 VPWR VGND sg13g2_decap_8
XFILLER_3_463 VPWR VGND sg13g2_decap_4
X_2070_ VPWR _1927_ net959 VGND sg13g2_inv_1
XFILLER_47_684 VPWR VGND sg13g2_decap_8
XFILLER_46_172 VPWR VGND sg13g2_decap_4
X_2972_ _1095_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ net636 VPWR VGND sg13g2_nand2_1
XFILLER_30_551 VPWR VGND sg13g2_decap_8
Xhold703 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] VPWR VGND net1022 sg13g2_dlygate4sd3_1
X_3524_ VGND VPWR _1913_ net585 _0308_ _1460_ sg13g2_a21oi_1
Xhold714 u_usb_cdc.sie_out_data\[3\] VPWR VGND net1033 sg13g2_dlygate4sd3_1
Xhold725 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[1\] VPWR VGND
+ net1044 sg13g2_dlygate4sd3_1
X_3455_ VGND VPWR net722 _1412_ _0285_ _1414_ sg13g2_a21oi_1
X_2406_ _0542_ _0634_ net744 _0636_ VPWR VGND sg13g2_nand3_1
X_3386_ net639 u_usb_cdc.sie_in_req _1371_ _1372_ VPWR VGND sg13g2_a21o_1
X_2337_ _0569_ net847 _0517_ VPWR VGND sg13g2_nand2_1
X_2268_ _0491_ _0483_ _0500_ VPWR VGND sg13g2_xor2_1
X_4007_ _2028_ _1009_ _1836_ _1840_ _1841_ VPWR VGND sg13g2_nor4_1
XFILLER_37_150 VPWR VGND sg13g2_fill_1
X_2199_ _0431_ VPWR _0432_ VGND net572 _2043_ sg13g2_o21ai_1
XFILLER_21_551 VPWR VGND sg13g2_fill_1
XFILLER_20_32 VPWR VGND sg13g2_fill_2
XFILLER_1_912 VPWR VGND sg13g2_decap_8
XFILLER_0_400 VPWR VGND sg13g2_decap_8
XFILLER_49_905 VPWR VGND sg13g2_decap_8
XFILLER_0_477 VPWR VGND sg13g2_decap_8
XFILLER_1_989 VPWR VGND sg13g2_decap_8
Xhold41 u_usb_cdc.u_sie.in_zlp_q\[1\] VPWR VGND net84 sg13g2_dlygate4sd3_1
Xhold30 _0104_ VPWR VGND net73 sg13g2_dlygate4sd3_1
XFILLER_21_1011 VPWR VGND sg13g2_decap_8
Xhold52 _0103_ VPWR VGND net95 sg13g2_dlygate4sd3_1
Xhold74 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[45\] VPWR VGND
+ net117 sg13g2_dlygate4sd3_1
Xhold63 _0098_ VPWR VGND net106 sg13g2_dlygate4sd3_1
Xhold85 _0210_ VPWR VGND net128 sg13g2_dlygate4sd3_1
Xhold96 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[69\] VPWR VGND
+ net139 sg13g2_dlygate4sd3_1
XFILLER_45_51 VPWR VGND sg13g2_fill_2
XFILLER_43_153 VPWR VGND sg13g2_fill_1
X_3240_ _1247_ VPWR _0237_ VGND _1155_ _1190_ sg13g2_o21ai_1
X_3171_ _1211_ net246 net609 VPWR VGND sg13g2_nand2_1
X_2122_ VPWR _1979_ net924 VGND sg13g2_inv_1
X_2053_ VPWR _1910_ net764 VGND sg13g2_inv_1
XFILLER_47_481 VPWR VGND sg13g2_decap_8
XFILLER_23_827 VPWR VGND sg13g2_decap_8
X_2955_ _1082_ VPWR _0116_ VGND net620 _1083_ sg13g2_o21ai_1
X_2886_ _1040_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net645 VPWR VGND sg13g2_nand2_1
Xhold511 _1809_ VPWR VGND net554 sg13g2_dlygate4sd3_1
Xhold500 u_usb_cdc.out_valid_o[0] VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold522 _0294_ VPWR VGND net565 sg13g2_dlygate4sd3_1
Xhold544 _0156_ VPWR VGND net863 sg13g2_dlygate4sd3_1
Xhold533 _0164_ VPWR VGND net852 sg13g2_dlygate4sd3_1
X_3507_ _1452_ net778 net775 VPWR VGND sg13g2_nand2_1
Xhold555 u_usb_cdc.u_ctrl_endp.req_q\[4\] VPWR VGND net874 sg13g2_dlygate4sd3_1
Xhold588 _0329_ VPWR VGND net907 sg13g2_dlygate4sd3_1
X_4487_ net733 VGND VPWR net47 u_usb_cdc.u_sie.u_phy_rx.dp_q\[0\] clknet_leaf_30_clk_regs
+ sg13g2_dfrbpq_1
Xhold577 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[12\] VPWR VGND net896 sg13g2_dlygate4sd3_1
Xhold566 net31 VPWR VGND net885 sg13g2_dlygate4sd3_1
X_3438_ net559 net582 _1405_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_9_clk_regs clknet_3_2__leaf_clk_regs clknet_leaf_9_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold599 _1803_ VPWR VGND net918 sg13g2_dlygate4sd3_1
X_3369_ net935 _1269_ _1360_ _0252_ VPWR VGND sg13g2_mux2_1
XFILLER_39_960 VPWR VGND sg13g2_decap_8
XFILLER_26_621 VPWR VGND sg13g2_decap_4
XFILLER_26_610 VPWR VGND sg13g2_fill_2
Xclkbuf_3_5__f_clk_regs clknet_0_clk_regs clknet_3_5__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_40_156 VPWR VGND sg13g2_fill_1
XFILLER_5_514 VPWR VGND sg13g2_fill_1
XFILLER_5_525 VPWR VGND sg13g2_fill_1
Xoutput31 net31 usb_dp_up_o VPWR VGND sg13g2_buf_1
XFILLER_1_720 VPWR VGND sg13g2_decap_8
Xoutput20 net20 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_49_702 VPWR VGND sg13g2_decap_8
XFILLER_0_274 VPWR VGND sg13g2_decap_8
XFILLER_1_797 VPWR VGND sg13g2_decap_8
XFILLER_49_779 VPWR VGND sg13g2_decap_8
XFILLER_45_974 VPWR VGND sg13g2_decap_8
XFILLER_31_101 VPWR VGND sg13g2_fill_2
XFILLER_20_819 VPWR VGND sg13g2_decap_8
X_2740_ _0930_ _0694_ _0744_ VPWR VGND sg13g2_nand2_1
XFILLER_12_392 VPWR VGND sg13g2_decap_4
X_2671_ _0876_ net841 net596 VPWR VGND sg13g2_nand2_1
X_4410_ net696 VGND VPWR _0338_ u_usb_cdc.u_sie.crc16_q\[15\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
X_4341_ net683 VGND VPWR _0269_ u_usb_cdc.addr\[1\] clknet_leaf_48_clk_regs sg13g2_dfrbpq_2
X_4272_ net654 VGND VPWR net181 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[34\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
XFILLER_28_1028 VPWR VGND sg13g2_fill_1
X_3223_ net758 net603 _1239_ VPWR VGND sg13g2_nor2_1
X_3154_ _1202_ net160 net607 VPWR VGND sg13g2_nand2_1
XFILLER_11_0 VPWR VGND sg13g2_fill_1
X_3085_ _1155_ net739 _1154_ VPWR VGND sg13g2_nand2_2
X_2105_ _1962_ net530 VPWR VGND sg13g2_inv_2
XFILLER_35_484 VPWR VGND sg13g2_fill_1
X_3987_ _1821_ VPWR _1822_ VGND _1921_ net709 sg13g2_o21ai_1
XFILLER_31_690 VPWR VGND sg13g2_fill_1
X_2938_ _1075_ VPWR _0106_ VGND net621 _1076_ sg13g2_o21ai_1
XFILLER_11_1010 VPWR VGND sg13g2_decap_8
X_2869_ net7 net1002 net646 _0080_ VPWR VGND sg13g2_mux2_1
Xhold330 _0229_ VPWR VGND net373 sg13g2_dlygate4sd3_1
Xhold341 _0413_ VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold352 _0033_ VPWR VGND net395 sg13g2_dlygate4sd3_1
Xhold385 u_usb_cdc.u_ctrl_endp.addr_dd\[2\] VPWR VGND net428 sg13g2_dlygate4sd3_1
Xhold374 _0217_ VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold363 u_usb_cdc.u_sie.in_toggle_q\[0\] VPWR VGND net406 sg13g2_dlygate4sd3_1
Xhold396 u_usb_cdc.u_sie.u_phy_tx.data_q\[2\] VPWR VGND net439 sg13g2_dlygate4sd3_1
Xfanout821 net825 net821 VPWR VGND sg13g2_buf_8
Xfanout832 net1046 net832 VPWR VGND sg13g2_buf_8
Xfanout843 net1026 net843 VPWR VGND sg13g2_buf_8
Xfanout810 net811 net810 VPWR VGND sg13g2_buf_8
XFILLER_26_53 VPWR VGND sg13g2_decap_8
XFILLER_27_996 VPWR VGND sg13g2_decap_8
XFILLER_42_966 VPWR VGND sg13g2_decap_8
XFILLER_26_484 VPWR VGND sg13g2_decap_8
XFILLER_13_178 VPWR VGND sg13g2_fill_2
XFILLER_6_801 VPWR VGND sg13g2_fill_1
XFILLER_10_841 VPWR VGND sg13g2_decap_8
XFILLER_10_874 VPWR VGND sg13g2_fill_1
XFILLER_5_344 VPWR VGND sg13g2_fill_2
XFILLER_1_594 VPWR VGND sg13g2_fill_1
XFILLER_1_583 VPWR VGND sg13g2_decap_8
XFILLER_1_572 VPWR VGND sg13g2_fill_2
XFILLER_49_576 VPWR VGND sg13g2_decap_8
XFILLER_17_484 VPWR VGND sg13g2_decap_8
X_3910_ net340 _1772_ _1775_ VPWR VGND sg13g2_and2_1
X_3841_ _1934_ _0450_ _0452_ _0481_ _1726_ VPWR VGND sg13g2_or4_1
XFILLER_20_605 VPWR VGND sg13g2_decap_4
XFILLER_32_498 VPWR VGND sg13g2_decap_4
XFILLER_20_649 VPWR VGND sg13g2_fill_1
X_3772_ VPWR VGND _1499_ net627 _1671_ net638 _1672_ _1669_ sg13g2_a221oi_1
X_2723_ _0919_ net393 _0918_ VPWR VGND sg13g2_nand2_1
X_2654_ _0865_ net766 _0864_ VPWR VGND sg13g2_nand2_1
X_2585_ _1942_ _0632_ _0636_ _0745_ _0808_ VPWR VGND sg13g2_nor4_1
X_4324_ net653 VGND VPWR net941 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[2\]
+ clknet_leaf_9_clk_regs sg13g2_dfrbpq_2
X_4255_ net655 VGND VPWR net442 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[17\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_3206_ VGND VPWR _1917_ net631 _0221_ _1229_ sg13g2_a21oi_1
X_4186_ net680 VGND VPWR net159 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[32\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
X_3137_ _1192_ net757 _1141_ VPWR VGND sg13g2_nand2_2
XFILLER_28_738 VPWR VGND sg13g2_fill_1
X_3068_ _1144_ VPWR _0168_ VGND net722 net635 sg13g2_o21ai_1
XFILLER_24_977 VPWR VGND sg13g2_decap_8
Xhold171 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[40\] VPWR
+ VGND net214 sg13g2_dlygate4sd3_1
Xhold160 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[8\] VPWR VGND
+ net203 sg13g2_dlygate4sd3_1
XFILLER_2_358 VPWR VGND sg13g2_decap_8
Xhold182 _0223_ VPWR VGND net225 sg13g2_dlygate4sd3_1
Xhold193 u_usb_cdc.u_sie.rx_data\[5\] VPWR VGND net236 sg13g2_dlygate4sd3_1
Xfanout651 net653 net651 VPWR VGND sg13g2_buf_8
Xfanout640 net641 net640 VPWR VGND sg13g2_buf_8
Xfanout684 net685 net684 VPWR VGND sg13g2_buf_8
Xfanout673 net674 net673 VPWR VGND sg13g2_buf_8
Xfanout662 net664 net662 VPWR VGND sg13g2_buf_8
Xfanout695 net704 net695 VPWR VGND sg13g2_buf_8
XFILLER_18_237 VPWR VGND sg13g2_fill_1
XFILLER_15_933 VPWR VGND sg13g2_fill_1
XFILLER_14_498 VPWR VGND sg13g2_decap_8
XFILLER_30_947 VPWR VGND sg13g2_decap_8
X_2370_ net752 _0600_ _0601_ VPWR VGND sg13g2_nor2_2
X_4040_ _1842_ VPWR _1870_ VGND u_usb_cdc.u_sie.u_phy_tx.data_q\[6\] _1835_ sg13g2_o21ai_1
Xclkbuf_leaf_23_clk_regs clknet_3_6__leaf_clk_regs clknet_leaf_23_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_21_936 VPWR VGND sg13g2_fill_1
X_3824_ _0357_ _1709_ _1711_ _1703_ _1934_ VPWR VGND sg13g2_a22oi_1
X_3755_ net776 _1514_ _1656_ VPWR VGND sg13g2_nor2b_1
X_2706_ _0883_ _0904_ _2042_ _0905_ VPWR VGND sg13g2_nand3_1
X_3686_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[19\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[27\]
+ net803 _1589_ VPWR VGND sg13g2_mux2_1
X_2637_ _0848_ u_usb_cdc.addr\[4\] u_usb_cdc.u_sie.addr_q\[4\] VPWR VGND sg13g2_xnor2_1
XFILLER_0_818 VPWR VGND sg13g2_decap_8
X_2568_ _0793_ _0643_ _0666_ VPWR VGND sg13g2_nand2_1
X_2499_ _0726_ net794 _0706_ VPWR VGND sg13g2_nand2_1
X_4307_ net650 VGND VPWR net227 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[69\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
X_4238_ net675 VGND VPWR net217 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[0\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
X_4169_ net678 VGND VPWR net106 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[15\]
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
XFILLER_28_568 VPWR VGND sg13g2_fill_2
XFILLER_23_284 VPWR VGND sg13g2_fill_1
XFILLER_47_866 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_546 VPWR VGND sg13g2_fill_1
XFILLER_19_557 VPWR VGND sg13g2_fill_2
XFILLER_34_505 VPWR VGND sg13g2_decap_8
XFILLER_46_365 VPWR VGND sg13g2_fill_2
XFILLER_46_376 VPWR VGND sg13g2_fill_1
XFILLER_14_284 VPWR VGND sg13g2_fill_1
XFILLER_30_755 VPWR VGND sg13g2_fill_2
XFILLER_31_1002 VPWR VGND sg13g2_decap_8
X_3540_ _1471_ net413 _1466_ VPWR VGND sg13g2_nand2_1
XFILLER_7_951 VPWR VGND sg13g2_decap_8
X_3471_ u_usb_cdc.sie_out_data\[2\] _1421_ _1426_ VPWR VGND sg13g2_nor2_1
X_2422_ _0652_ net792 net785 VPWR VGND sg13g2_nand2_1
X_2353_ net327 net321 net376 _0584_ VPWR VGND sg13g2_nand3_1
X_2284_ _0516_ net710 VPWR VGND net768 sg13g2_nand2b_2
X_4023_ _1852_ _1853_ _0926_ _1855_ VPWR VGND _1854_ sg13g2_nand4_1
XFILLER_25_549 VPWR VGND sg13g2_decap_8
XFILLER_33_582 VPWR VGND sg13g2_fill_2
XFILLER_21_755 VPWR VGND sg13g2_fill_2
X_3807_ net592 _1692_ net992 _1699_ VPWR VGND sg13g2_nand3_1
X_3738_ net804 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[5\] _1639_
+ VPWR VGND sg13g2_nor2b_1
X_3669_ VPWR VGND _1569_ _1572_ _1567_ _1500_ _1573_ _1564_ sg13g2_a221oi_1
XFILLER_47_1020 VPWR VGND sg13g2_decap_8
XFILLER_48_619 VPWR VGND sg13g2_decap_8
XFILLER_47_129 VPWR VGND sg13g2_fill_2
XFILLER_29_877 VPWR VGND sg13g2_decap_4
XFILLER_34_42 VPWR VGND sg13g2_fill_2
XFILLER_7_236 VPWR VGND sg13g2_fill_2
XFILLER_3_420 VPWR VGND sg13g2_fill_2
XFILLER_38_118 VPWR VGND sg13g2_fill_1
XFILLER_47_663 VPWR VGND sg13g2_decap_8
X_2971_ _1094_ net177 _1079_ VPWR VGND sg13g2_nand2_1
XFILLER_43_891 VPWR VGND sg13g2_decap_8
XFILLER_15_582 VPWR VGND sg13g2_decap_4
XFILLER_30_596 VPWR VGND sg13g2_fill_1
Xhold704 _0064_ VPWR VGND net1023 sg13g2_dlygate4sd3_1
Xhold726 u_usb_cdc.sie_out_data\[2\] VPWR VGND net1045 sg13g2_dlygate4sd3_1
X_3523_ net385 net585 _1460_ VPWR VGND sg13g2_nor2_1
Xhold715 u_usb_cdc.sie_in_req VPWR VGND net1034 sg13g2_dlygate4sd3_1
X_3454_ net953 _1412_ _1414_ VPWR VGND sg13g2_nor2_1
X_2405_ _0635_ _0633_ VPWR VGND net779 sg13g2_nand2b_2
X_3385_ net809 net801 net797 _1371_ VGND VPWR _1924_ sg13g2_nor4_2
X_2336_ VPWR VGND net84 _0565_ net638 net164 _0568_ net640 sg13g2_a221oi_1
X_2267_ _0499_ u_usb_cdc.u_sie.crc16_q\[1\] _0484_ VPWR VGND sg13g2_xnor2_1
X_4006_ VGND VPWR _0926_ _1839_ _1840_ _1834_ sg13g2_a21oi_1
X_2198_ _0431_ net990 net707 VPWR VGND sg13g2_nand2_1
Xclkbuf_3_4__f_clk_regs clknet_0_clk_regs clknet_3_4__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_1_968 VPWR VGND sg13g2_decap_8
XFILLER_0_456 VPWR VGND sg13g2_decap_8
Xhold31 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[42\] VPWR VGND
+ net74 sg13g2_dlygate4sd3_1
Xhold20 _0123_ VPWR VGND net63 sg13g2_dlygate4sd3_1
Xhold64 u_usb_cdc.u_sie.out_eop_q VPWR VGND net107 sg13g2_dlygate4sd3_1
Xhold42 _0425_ VPWR VGND net85 sg13g2_dlygate4sd3_1
Xhold53 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[47\] VPWR VGND
+ net96 sg13g2_dlygate4sd3_1
Xhold86 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[65\] VPWR VGND
+ net129 sg13g2_dlygate4sd3_1
Xhold75 _0128_ VPWR VGND net118 sg13g2_dlygate4sd3_1
Xhold97 _0152_ VPWR VGND net140 sg13g2_dlygate4sd3_1
XFILLER_12_563 VPWR VGND sg13g2_decap_4
XFILLER_12_585 VPWR VGND sg13g2_fill_2
XFILLER_3_294 VPWR VGND sg13g2_fill_1
X_3170_ _1210_ VPWR _0204_ VGND _1188_ net608 sg13g2_o21ai_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_13_4 VPWR VGND sg13g2_fill_1
X_2121_ _1978_ net929 VPWR VGND sg13g2_inv_2
X_2052_ VPWR _1909_ net299 VGND sg13g2_inv_1
XFILLER_48_983 VPWR VGND sg13g2_decap_8
X_2954_ _1083_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2885_ net833 net834 _1039_ VPWR VGND sg13g2_nor2b_2
Xhold501 _0042_ VPWR VGND net544 sg13g2_dlygate4sd3_1
Xhold512 _0396_ VPWR VGND net555 sg13g2_dlygate4sd3_1
Xhold523 u_usb_cdc.u_ctrl_endp.addr_dd\[4\] VPWR VGND net566 sg13g2_dlygate4sd3_1
Xhold545 u_usb_cdc.u_ctrl_endp.max_length_q\[2\] VPWR VGND net864 sg13g2_dlygate4sd3_1
X_3506_ _1451_ net774 _1437_ VPWR VGND sg13g2_nand2_1
Xhold534 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] VPWR VGND net853 sg13g2_dlygate4sd3_1
Xhold556 _0005_ VPWR VGND net875 sg13g2_dlygate4sd3_1
Xhold578 u_usb_cdc.addr\[4\] VPWR VGND net897 sg13g2_dlygate4sd3_1
Xhold567 _1820_ VPWR VGND net886 sg13g2_dlygate4sd3_1
X_4486_ net735 VGND VPWR net887 net31 clknet_leaf_26_clk_regs sg13g2_dfrbpq_2
XFILLER_44_1012 VPWR VGND sg13g2_decap_8
X_3437_ VGND VPWR _1913_ net581 _0277_ _1404_ sg13g2_a21oi_1
Xhold589 u_usb_cdc.u_ctrl_endp.max_length_q\[5\] VPWR VGND net908 sg13g2_dlygate4sd3_1
X_3368_ _1361_ VPWR _0251_ VGND _1984_ _1360_ sg13g2_o21ai_1
X_2319_ u_usb_cdc.u_ctrl_endp.state_q\[1\] u_usb_cdc.ctrl_stall u_usb_cdc.u_ctrl_endp.state_q\[5\]
+ _0550_ _0551_ VPWR VGND sg13g2_or4_1
X_3299_ _1299_ VPWR _1300_ VGND net822 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[17\]
+ sg13g2_o21ai_1
XFILLER_14_806 VPWR VGND sg13g2_fill_2
XFILLER_26_677 VPWR VGND sg13g2_fill_1
XFILLER_15_55 VPWR VGND sg13g2_fill_2
XFILLER_22_894 VPWR VGND sg13g2_fill_2
XFILLER_40_179 VPWR VGND sg13g2_fill_1
Xoutput21 net21 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_1_776 VPWR VGND sg13g2_decap_8
XFILLER_0_253 VPWR VGND sg13g2_decap_8
XFILLER_0_242 VPWR VGND sg13g2_fill_1
XFILLER_49_758 VPWR VGND sg13g2_decap_8
XFILLER_45_953 VPWR VGND sg13g2_decap_8
XFILLER_16_121 VPWR VGND sg13g2_fill_1
XFILLER_32_603 VPWR VGND sg13g2_decap_8
XFILLER_13_850 VPWR VGND sg13g2_fill_1
X_2670_ net1027 VPWR _0026_ VGND _0572_ _0590_ sg13g2_o21ai_1
Xclkbuf_leaf_48_clk_regs clknet_3_4__leaf_clk_regs clknet_leaf_48_clk_regs VPWR VGND
+ sg13g2_buf_8
X_4340_ net684 VGND VPWR _0268_ u_usb_cdc.addr\[0\] clknet_leaf_44_clk_regs sg13g2_dfrbpq_2
XFILLER_28_1007 VPWR VGND sg13g2_decap_8
X_4271_ net655 VGND VPWR net144 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[33\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_3222_ _1238_ VPWR _0228_ VGND _1914_ net603 sg13g2_o21ai_1
X_3153_ VGND VPWR _1999_ net605 _0196_ _1201_ sg13g2_a21oi_1
X_2104_ VPWR _1961_ net915 VGND sg13g2_inv_1
X_3084_ net827 _1153_ _1154_ VPWR VGND sg13g2_nor2_2
XFILLER_48_780 VPWR VGND sg13g2_decap_8
XFILLER_36_986 VPWR VGND sg13g2_decap_8
XFILLER_23_647 VPWR VGND sg13g2_decap_4
X_3986_ _1821_ _0433_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] _2027_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_2937_ _1076_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ _1059_ VPWR VGND sg13g2_nand2_1
X_2868_ net6 net1000 net646 _0079_ VPWR VGND sg13g2_mux2_1
X_2799_ net750 VPWR _0975_ VGND net839 _0974_ sg13g2_o21ai_1
Xhold320 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[3\] VPWR VGND
+ net363 sg13g2_dlygate4sd3_1
Xhold342 u_usb_cdc.u_sie.addr_q\[2\] VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold353 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[55\] VPWR
+ VGND net396 sg13g2_dlygate4sd3_1
Xhold331 u_usb_cdc.u_sie.u_phy_rx.se0_q VPWR VGND net374 sg13g2_dlygate4sd3_1
Xhold375 u_usb_cdc.u_ctrl_endp.endp_q\[0\] VPWR VGND net418 sg13g2_dlygate4sd3_1
Xhold386 _0277_ VPWR VGND net429 sg13g2_dlygate4sd3_1
XFILLER_7_9 VPWR VGND sg13g2_fill_1
Xhold364 _0069_ VPWR VGND net407 sg13g2_dlygate4sd3_1
X_4469_ net734 VGND VPWR net307 u_usb_cdc.u_sie.u_phy_rx.rx_err_q clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_1
Xfanout800 net802 net800 VPWR VGND sg13g2_buf_8
Xhold397 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[17\] VPWR
+ VGND net440 sg13g2_dlygate4sd3_1
Xfanout822 net823 net822 VPWR VGND sg13g2_buf_1
Xfanout833 net1044 net833 VPWR VGND sg13g2_buf_8
Xfanout811 net1038 net811 VPWR VGND sg13g2_buf_8
Xfanout844 net921 net844 VPWR VGND sg13g2_buf_8
XFILLER_46_739 VPWR VGND sg13g2_decap_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_27_975 VPWR VGND sg13g2_decap_8
XFILLER_42_945 VPWR VGND sg13g2_decap_8
XFILLER_13_157 VPWR VGND sg13g2_fill_2
XFILLER_42_20 VPWR VGND sg13g2_fill_2
XFILLER_9_128 VPWR VGND sg13g2_fill_2
XFILLER_42_31 VPWR VGND sg13g2_decap_4
XFILLER_49_555 VPWR VGND sg13g2_decap_8
XFILLER_45_794 VPWR VGND sg13g2_decap_8
X_3840_ net752 net717 _0436_ _0950_ _1725_ VPWR VGND sg13g2_nor4_1
X_3771_ _1652_ VPWR _1671_ VGND _1630_ _1670_ sg13g2_o21ai_1
XFILLER_34_1022 VPWR VGND sg13g2_decap_8
X_2722_ net391 net457 net744 _0918_ VPWR VGND sg13g2_nand3_1
X_2653_ _0854_ _0857_ _0863_ _0864_ VPWR VGND sg13g2_nor3_1
X_2584_ _0664_ _0699_ _0651_ _0807_ VPWR VGND _0806_ sg13g2_nand4_1
X_4323_ net653 VGND VPWR net936 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[1\]
+ clknet_leaf_9_clk_regs sg13g2_dfrbpq_2
X_4254_ net656 VGND VPWR net399 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[16\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
XFILLER_41_1026 VPWR VGND sg13g2_fill_2
X_3205_ net426 net631 _1229_ VPWR VGND sg13g2_nor2_1
X_4185_ net678 VGND VPWR net510 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[31\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
X_3136_ net333 net633 _1191_ VPWR VGND sg13g2_nor2_1
XFILLER_27_216 VPWR VGND sg13g2_fill_1
X_3067_ _1144_ net252 _1142_ VPWR VGND sg13g2_nand2_1
X_3969_ _1813_ net187 net614 VPWR VGND sg13g2_nand2_1
XFILLER_2_337 VPWR VGND sg13g2_decap_8
Xhold150 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[9\] VPWR VGND
+ net193 sg13g2_dlygate4sd3_1
Xhold161 _0175_ VPWR VGND net204 sg13g2_dlygate4sd3_1
Xhold172 _0207_ VPWR VGND net215 sg13g2_dlygate4sd3_1
Xhold183 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[69\] VPWR
+ VGND net226 sg13g2_dlygate4sd3_1
Xhold194 _0406_ VPWR VGND net237 sg13g2_dlygate4sd3_1
Xfanout630 net631 net630 VPWR VGND sg13g2_buf_8
Xfanout641 _0515_ net641 VPWR VGND sg13g2_buf_8
Xfanout685 net690 net685 VPWR VGND sg13g2_buf_8
Xfanout674 net675 net674 VPWR VGND sg13g2_buf_8
Xfanout652 net653 net652 VPWR VGND sg13g2_buf_8
XFILLER_19_706 VPWR VGND sg13g2_fill_1
Xfanout663 net665 net663 VPWR VGND sg13g2_buf_8
Xfanout696 net704 net696 VPWR VGND sg13g2_buf_2
XFILLER_19_717 VPWR VGND sg13g2_fill_1
XFILLER_18_1017 VPWR VGND sg13g2_decap_8
XFILLER_42_764 VPWR VGND sg13g2_fill_2
XFILLER_30_926 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_4
XFILLER_1_381 VPWR VGND sg13g2_decap_8
XFILLER_49_330 VPWR VGND sg13g2_fill_1
XFILLER_37_536 VPWR VGND sg13g2_fill_1
XFILLER_17_282 VPWR VGND sg13g2_fill_2
XFILLER_33_753 VPWR VGND sg13g2_fill_2
X_3823_ VGND VPWR net765 _1710_ _1711_ _1703_ sg13g2_a21oi_1
X_3754_ net773 _0544_ _1654_ _1655_ VPWR VGND sg13g2_nor3_1
X_2705_ VPWR _0904_ _0903_ VGND sg13g2_inv_1
X_3685_ VGND VPWR net803 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[11\]
+ _1588_ _1587_ sg13g2_a21oi_1
X_2636_ _0847_ u_usb_cdc.addr\[3\] u_usb_cdc.u_sie.addr_q\[3\] VPWR VGND sg13g2_xnor2_1
X_2567_ _0610_ _0615_ net591 _0792_ VPWR VGND sg13g2_nor3_1
X_2498_ _0725_ _0693_ _0711_ _0724_ VPWR VGND sg13g2_and3_1
X_4306_ net649 VGND VPWR _0235_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[68\]
+ clknet_3_0__leaf_clk_regs sg13g2_dfrbpq_1
X_4237_ net681 VGND VPWR net364 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[3\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_2
X_4168_ net662 VGND VPWR net221 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[14\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_4099_ net690 VGND VPWR net514 u_usb_cdc.u_ctrl_endp.req_q\[5\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
X_3119_ _1180_ net762 _1141_ VPWR VGND sg13g2_nand2_2
XFILLER_16_709 VPWR VGND sg13g2_fill_1
XFILLER_24_742 VPWR VGND sg13g2_decap_4
XFILLER_12_915 VPWR VGND sg13g2_fill_2
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_48_85 VPWR VGND sg13g2_fill_2
XFILLER_47_845 VPWR VGND sg13g2_decap_8
X_3470_ net864 net576 _1425_ VPWR VGND sg13g2_nor2_1
X_2421_ _0651_ net588 _0643_ _0650_ VPWR VGND sg13g2_and3_1
X_2352_ _0574_ net988 _0583_ _0063_ VPWR VGND sg13g2_nor3_1
X_2283_ net769 _2015_ _0515_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_812 VPWR VGND sg13g2_fill_2
X_4022_ _1854_ _2027_ net292 VPWR VGND sg13g2_nand2b_1
XFILLER_18_591 VPWR VGND sg13g2_fill_1
Xclkbuf_3_3__f_clk_regs clknet_0_clk_regs clknet_3_3__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_21_723 VPWR VGND sg13g2_decap_8
XFILLER_21_712 VPWR VGND sg13g2_fill_2
XFILLER_20_200 VPWR VGND sg13g2_fill_2
X_3806_ _1698_ VPWR _0352_ VGND _1914_ net600 sg13g2_o21ai_1
X_3737_ _1638_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[69\] net628
+ VPWR VGND sg13g2_nand2_1
X_3668_ _1571_ net773 _1513_ _1572_ VPWR VGND sg13g2_a21o_1
X_3599_ _1500_ VPWR _1505_ VGND _1502_ _1504_ sg13g2_o21ai_1
X_2619_ _0833_ VPWR _0015_ VGND _0820_ _0825_ sg13g2_o21ai_1
XFILLER_24_594 VPWR VGND sg13g2_fill_1
XFILLER_24_583 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_4_988 VPWR VGND sg13g2_decap_8
XFILLER_47_642 VPWR VGND sg13g2_decap_8
XFILLER_15_550 VPWR VGND sg13g2_fill_1
X_2970_ _1092_ VPWR _0121_ VGND net621 _1093_ sg13g2_o21ai_1
XFILLER_30_586 VPWR VGND sg13g2_fill_2
Xhold705 u_usb_cdc.sie_out_data\[6\] VPWR VGND net1024 sg13g2_dlygate4sd3_1
X_3522_ VGND VPWR net721 net586 _0307_ _1459_ sg13g2_a21oi_1
Xhold727 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[0\] VPWR
+ VGND net1046 sg13g2_dlygate4sd3_1
Xhold716 u_usb_cdc.u_sie.phy_state_q\[4\] VPWR VGND net1035 sg13g2_dlygate4sd3_1
X_3453_ VGND VPWR net724 _1412_ _0284_ _1413_ sg13g2_a21oi_1
X_2404_ net779 net772 _0546_ _0634_ VPWR VGND sg13g2_nor3_2
X_3384_ net931 net639 net1034 _1370_ VPWR VGND sg13g2_nand3_1
X_2335_ net769 _2015_ _0567_ VPWR VGND sg13g2_and2_1
X_2266_ _0498_ _1962_ _0485_ VPWR VGND sg13g2_xnor2_1
X_2197_ _0430_ _0429_ net990 VPWR VGND sg13g2_nand2b_1
X_4005_ _1837_ _1838_ _2018_ _1839_ VPWR VGND sg13g2_nand3_1
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_38_686 VPWR VGND sg13g2_decap_4
XFILLER_38_1009 VPWR VGND sg13g2_decap_8
XFILLER_26_859 VPWR VGND sg13g2_fill_2
XFILLER_21_542 VPWR VGND sg13g2_decap_8
XFILLER_4_218 VPWR VGND sg13g2_fill_2
XFILLER_0_435 VPWR VGND sg13g2_decap_8
XFILLER_1_947 VPWR VGND sg13g2_decap_8
Xhold10 u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[0\] VPWR VGND net53 sg13g2_dlygate4sd3_1
XFILLER_29_32 VPWR VGND sg13g2_decap_4
Xhold32 _0125_ VPWR VGND net75 sg13g2_dlygate4sd3_1
Xhold21 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[41\] VPWR VGND
+ net64 sg13g2_dlygate4sd3_1
Xhold43 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[51\] VPWR VGND
+ net86 sg13g2_dlygate4sd3_1
Xhold65 _0360_ VPWR VGND net108 sg13g2_dlygate4sd3_1
Xhold54 _0130_ VPWR VGND net97 sg13g2_dlygate4sd3_1
Xhold87 _0232_ VPWR VGND net130 sg13g2_dlygate4sd3_1
Xhold98 _0050_ VPWR VGND net141 sg13g2_dlygate4sd3_1
XFILLER_29_642 VPWR VGND sg13g2_decap_8
Xhold76 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[12\] VPWR VGND
+ net119 sg13g2_dlygate4sd3_1
XFILLER_45_31 VPWR VGND sg13g2_fill_1
XFILLER_44_601 VPWR VGND sg13g2_fill_1
XFILLER_45_53 VPWR VGND sg13g2_fill_1
XFILLER_43_166 VPWR VGND sg13g2_fill_1
XFILLER_8_546 VPWR VGND sg13g2_decap_4
XFILLER_6_1007 VPWR VGND sg13g2_decap_8
X_2120_ VPWR _1977_ u_usb_cdc.u_sie.u_phy_rx.state_q\[2\] VGND sg13g2_inv_1
XFILLER_48_962 VPWR VGND sg13g2_decap_8
X_2051_ VPWR _1908_ net481 VGND sg13g2_inv_1
XFILLER_47_450 VPWR VGND sg13g2_decap_8
XFILLER_34_144 VPWR VGND sg13g2_fill_1
XFILLER_37_1020 VPWR VGND sg13g2_decap_8
X_2953_ _1082_ net218 _1079_ VPWR VGND sg13g2_nand2_1
X_2884_ _1038_ net82 _1037_ VPWR VGND sg13g2_nand2_1
Xhold502 u_usb_cdc.u_ctrl_endp.endp_q\[2\] VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold524 u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[1\] VPWR VGND net567 sg13g2_dlygate4sd3_1
Xhold513 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\] VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold535 u_usb_cdc.u_sie.crc16_q\[2\] VPWR VGND net854 sg13g2_dlygate4sd3_1
X_3505_ _1448_ VPWR _0299_ VGND _1439_ _1450_ sg13g2_o21ai_1
X_4485_ net737 VGND VPWR _0047_ u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[1\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_1
Xhold579 u_usb_cdc.u_ctrl_endp.max_length_q\[3\] VPWR VGND net898 sg13g2_dlygate4sd3_1
Xhold546 _0290_ VPWR VGND net865 sg13g2_dlygate4sd3_1
Xhold557 u_usb_cdc.u_sie.rx_err VPWR VGND net876 sg13g2_dlygate4sd3_1
Xhold568 _0409_ VPWR VGND net887 sg13g2_dlygate4sd3_1
X_3436_ net428 net581 _1404_ VPWR VGND sg13g2_nor2_1
X_3367_ _1361_ _1266_ _1360_ VPWR VGND sg13g2_nand2_1
X_2318_ _0550_ net541 u_usb_cdc.u_ctrl_endp.state_q\[7\] VPWR VGND sg13g2_nand2b_1
X_3298_ _1299_ net822 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[25\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_39_995 VPWR VGND sg13g2_decap_8
X_2249_ _0481_ _0478_ _0441_ VPWR VGND sg13g2_nand2b_1
XFILLER_15_45 VPWR VGND sg13g2_fill_1
XFILLER_41_626 VPWR VGND sg13g2_decap_4
XFILLER_31_44 VPWR VGND sg13g2_decap_4
Xoutput22 net22 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_755 VPWR VGND sg13g2_decap_8
XFILLER_0_232 VPWR VGND sg13g2_fill_2
XFILLER_49_737 VPWR VGND sg13g2_decap_8
XFILLER_45_932 VPWR VGND sg13g2_decap_8
XFILLER_16_188 VPWR VGND sg13g2_fill_2
XFILLER_31_103 VPWR VGND sg13g2_fill_1
XFILLER_32_637 VPWR VGND sg13g2_decap_8
XFILLER_40_670 VPWR VGND sg13g2_decap_8
X_4270_ net658 VGND VPWR net258 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[32\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
X_3221_ _1238_ net323 net604 VPWR VGND sg13g2_nand2_1
X_3152_ u_usb_cdc.sie_out_data\[5\] net605 _1201_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_17_clk_regs clknet_3_3__leaf_clk_regs clknet_leaf_17_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2103_ VPWR _1960_ u_usb_cdc.u_sie.data_q\[6\] VGND sg13g2_inv_1
X_3083_ VGND VPWR _1153_ net829 net830 sg13g2_or2_1
XFILLER_22_103 VPWR VGND sg13g2_fill_2
XFILLER_22_125 VPWR VGND sg13g2_fill_2
X_3985_ VGND VPWR net748 _0921_ _0409_ net886 sg13g2_a21oi_1
X_2936_ _1075_ net121 _1060_ VPWR VGND sg13g2_nand2_1
X_2867_ net5 net996 net646 _0078_ VPWR VGND sg13g2_mux2_1
X_2798_ net767 _0973_ _0974_ VPWR VGND sg13g2_nor2_1
Xhold310 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[15\] VPWR VGND net353 sg13g2_dlygate4sd3_1
Xhold343 _0308_ VPWR VGND net386 sg13g2_dlygate4sd3_1
Xhold321 _0166_ VPWR VGND net364 sg13g2_dlygate4sd3_1
Xhold332 _0421_ VPWR VGND net375 sg13g2_dlygate4sd3_1
Xhold365 u_usb_cdc.u_sie.addr_q\[4\] VPWR VGND net408 sg13g2_dlygate4sd3_1
Xhold354 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[16\] VPWR
+ VGND net397 sg13g2_dlygate4sd3_1
Xhold387 u_usb_cdc.u_sie.delay_cnt_q\[1\] VPWR VGND net430 sg13g2_dlygate4sd3_1
X_4468_ net732 VGND VPWR _0395_ u_usb_cdc.u_sie.rx_valid clknet_leaf_32_clk_regs sg13g2_dfrbpq_1
Xhold376 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[2\] VPWR VGND
+ net419 sg13g2_dlygate4sd3_1
Xfanout823 net825 net823 VPWR VGND sg13g2_buf_8
Xhold398 _1179_ VPWR VGND net441 sg13g2_dlygate4sd3_1
Xfanout812 net813 net812 VPWR VGND sg13g2_buf_8
Xfanout801 net802 net801 VPWR VGND sg13g2_buf_8
X_3419_ u_usb_cdc.u_ctrl_endp.req_q\[7\] net849 _1396_ VPWR VGND sg13g2_nor2b_1
Xfanout834 net977 net834 VPWR VGND sg13g2_buf_8
X_4399_ net700 VGND VPWR _0327_ u_usb_cdc.u_sie.crc16_q\[4\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
Xfanout845 net846 net845 VPWR VGND sg13g2_buf_8
XFILLER_46_718 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_45_239 VPWR VGND sg13g2_decap_8
XFILLER_42_924 VPWR VGND sg13g2_decap_8
XFILLER_13_114 VPWR VGND sg13g2_fill_1
XFILLER_41_423 VPWR VGND sg13g2_decap_4
XFILLER_10_854 VPWR VGND sg13g2_decap_8
XFILLER_5_346 VPWR VGND sg13g2_fill_1
XFILLER_49_534 VPWR VGND sg13g2_decap_8
XFILLER_45_773 VPWR VGND sg13g2_decap_8
XFILLER_33_946 VPWR VGND sg13g2_fill_2
X_3770_ _0537_ VPWR _1670_ VGND net773 _0536_ sg13g2_o21ai_1
XFILLER_20_629 VPWR VGND sg13g2_fill_1
XFILLER_34_1001 VPWR VGND sg13g2_decap_8
X_2721_ _0917_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] _0916_ VPWR VGND sg13g2_nand2_1
XFILLER_9_696 VPWR VGND sg13g2_fill_1
X_2652_ _0863_ net767 _0862_ VPWR VGND sg13g2_nand2_1
X_2583_ _0637_ _0641_ _0667_ _0806_ VPWR VGND sg13g2_nor3_1
X_4322_ net652 VGND VPWR net1004 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[0\]
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
X_4253_ net657 VGND VPWR net116 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[15\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_3204_ VGND VPWR _1914_ net630 _0220_ _1228_ sg13g2_a21oi_1
XFILLER_41_1005 VPWR VGND sg13g2_decap_8
X_4184_ net664 VGND VPWR net571 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[30\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
X_3135_ VGND VPWR net632 _1190_ _0189_ _1189_ sg13g2_a21oi_1
X_3066_ _1143_ VPWR _0167_ VGND net723 net634 sg13g2_o21ai_1
X_3968_ _0988_ VPWR _0400_ VGND _1918_ net742 sg13g2_o21ai_1
X_2919_ _1064_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net644 VPWR VGND sg13g2_nand2_1
X_3899_ _1747_ _1765_ _1766_ _1767_ VPWR VGND sg13g2_nor3_1
Xhold140 _0101_ VPWR VGND net183 sg13g2_dlygate4sd3_1
Xhold151 _0092_ VPWR VGND net194 sg13g2_dlygate4sd3_1
Xhold162 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[36\] VPWR VGND
+ net205 sg13g2_dlygate4sd3_1
Xhold184 _0236_ VPWR VGND net227 sg13g2_dlygate4sd3_1
Xhold173 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[0\] VPWR VGND
+ net216 sg13g2_dlygate4sd3_1
Xhold195 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[22\] VPWR VGND
+ net238 sg13g2_dlygate4sd3_1
Xfanout631 _1222_ net631 VPWR VGND sg13g2_buf_8
Xfanout642 net643 net642 VPWR VGND sg13g2_buf_8
Xfanout620 net621 net620 VPWR VGND sg13g2_buf_8
Xfanout653 net671 net653 VPWR VGND sg13g2_buf_8
Xfanout675 net682 net675 VPWR VGND sg13g2_buf_8
Xfanout664 net665 net664 VPWR VGND sg13g2_buf_2
Xfanout686 net690 net686 VPWR VGND sg13g2_buf_8
XFILLER_19_729 VPWR VGND sg13g2_decap_8
Xfanout697 net699 net697 VPWR VGND sg13g2_buf_8
XFILLER_2_1010 VPWR VGND sg13g2_decap_8
XFILLER_37_43 VPWR VGND sg13g2_decap_4
XFILLER_42_732 VPWR VGND sg13g2_fill_1
XFILLER_30_905 VPWR VGND sg13g2_fill_2
XFILLER_10_651 VPWR VGND sg13g2_fill_1
XFILLER_6_633 VPWR VGND sg13g2_fill_2
XFILLER_5_165 VPWR VGND sg13g2_fill_2
XFILLER_1_360 VPWR VGND sg13g2_decap_8
XFILLER_18_762 VPWR VGND sg13g2_fill_2
Xclkbuf_3_2__f_clk_regs clknet_0_clk_regs clknet_3_2__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_32_220 VPWR VGND sg13g2_fill_1
XFILLER_33_765 VPWR VGND sg13g2_decap_4
X_3822_ _0862_ _1701_ _1710_ VPWR VGND sg13g2_and2_1
X_3753_ net780 _0543_ _0761_ _1503_ _1654_ VPWR VGND sg13g2_and4_1
X_2704_ _2038_ _0884_ net1007 _0903_ VPWR VGND sg13g2_nand3_1
X_3684_ net803 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[3\] _1587_
+ VPWR VGND sg13g2_nor2b_1
X_2635_ _0846_ u_usb_cdc.addr\[5\] u_usb_cdc.u_sie.addr_q\[5\] VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_32_clk_regs clknet_3_7__leaf_clk_regs clknet_leaf_32_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2566_ _0790_ VPWR _0006_ VGND _0708_ _0791_ sg13g2_o21ai_1
X_4305_ net649 VGND VPWR net192 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[67\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
X_2497_ _0724_ _0723_ _0459_ VPWR VGND sg13g2_nand2b_1
X_4236_ net679 VGND VPWR net420 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[2\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
X_4167_ net662 VGND VPWR net132 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[13\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
X_3118_ net440 net633 _1179_ VPWR VGND sg13g2_nor2_1
X_4098_ net689 VGND VPWR net875 u_usb_cdc.u_ctrl_endp.req_q\[4\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_2
X_3049_ _1028_ net1025 _1032_ _0161_ VPWR VGND sg13g2_mux2_1
XFILLER_24_776 VPWR VGND sg13g2_decap_8
XFILLER_24_787 VPWR VGND sg13g2_fill_1
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_47_824 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_46_367 VPWR VGND sg13g2_fill_1
XFILLER_7_986 VPWR VGND sg13g2_decap_8
X_2420_ _0611_ _0616_ _0630_ _0649_ _0650_ VPWR VGND sg13g2_or4_1
X_2351_ VPWR _0583_ _0582_ VGND sg13g2_inv_1
XFILLER_9_1016 VPWR VGND sg13g2_decap_8
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
X_2282_ net768 u_usb_cdc.endp\[1\] _0514_ VPWR VGND sg13g2_nor2_1
X_4021_ _1853_ _1979_ _2028_ VPWR VGND sg13g2_nand2_1
XFILLER_38_857 VPWR VGND sg13g2_fill_2
XFILLER_46_890 VPWR VGND sg13g2_decap_8
XFILLER_21_735 VPWR VGND sg13g2_fill_1
X_3805_ net592 _1692_ net989 _1698_ VPWR VGND sg13g2_nand3_1
XFILLER_20_256 VPWR VGND sg13g2_fill_2
X_3736_ _1637_ net989 net597 VPWR VGND sg13g2_nand2_1
X_3667_ VGND VPWR _0647_ _1441_ _1571_ _1570_ sg13g2_a21oi_1
X_3598_ _1504_ _1503_ _0544_ VPWR VGND sg13g2_nand2b_1
X_2618_ _0833_ net471 net591 VPWR VGND sg13g2_nand2_1
X_2549_ _0775_ _0648_ _0776_ VPWR VGND sg13g2_nor2b_1
X_4219_ net667 VGND VPWR net201 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[65\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
XFILLER_18_45 VPWR VGND sg13g2_fill_2
XFILLER_34_44 VPWR VGND sg13g2_fill_1
XFILLER_12_757 VPWR VGND sg13g2_decap_8
XFILLER_12_768 VPWR VGND sg13g2_fill_1
XFILLER_7_238 VPWR VGND sg13g2_fill_1
XFILLER_4_967 VPWR VGND sg13g2_decap_8
XFILLER_47_698 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_decap_8
X_3521_ net449 net586 _1459_ VPWR VGND sg13g2_nor2_1
XFILLER_6_271 VPWR VGND sg13g2_fill_2
Xhold728 u_usb_cdc.u_sie.phy_state_q\[1\] VPWR VGND net1047 sg13g2_dlygate4sd3_1
Xhold717 _0879_ VPWR VGND net1036 sg13g2_dlygate4sd3_1
Xhold706 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\] VPWR VGND
+ net1025 sg13g2_dlygate4sd3_1
X_3452_ net880 _1412_ _1413_ VPWR VGND sg13g2_nor2_1
X_2403_ net772 _0546_ _0633_ VPWR VGND sg13g2_nor2_2
X_3383_ _1369_ _1128_ _1134_ VPWR VGND sg13g2_nand2_2
X_2334_ u_usb_cdc.endp\[1\] net768 _0566_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
X_2265_ _0497_ _0490_ _0495_ VPWR VGND sg13g2_xnor2_1
X_2196_ _0429_ _2033_ _2031_ VPWR VGND sg13g2_nand2b_1
X_4004_ _1838_ _1954_ net845 u_usb_cdc.u_sie.pid_q\[1\] net836 VPWR VGND sg13g2_a22oi_1
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_41_808 VPWR VGND sg13g2_decap_4
XFILLER_14_1021 VPWR VGND sg13g2_decap_8
XFILLER_4_208 VPWR VGND sg13g2_fill_2
X_3719_ net798 _1619_ _1620_ _1621_ VPWR VGND sg13g2_nor3_1
XFILLER_20_68 VPWR VGND sg13g2_fill_1
XFILLER_1_926 VPWR VGND sg13g2_decap_8
XFILLER_0_414 VPWR VGND sg13g2_decap_8
XFILLER_29_11 VPWR VGND sg13g2_decap_8
Xhold11 _0046_ VPWR VGND net54 sg13g2_dlygate4sd3_1
XFILLER_49_919 VPWR VGND sg13g2_decap_8
Xhold22 _0124_ VPWR VGND net65 sg13g2_dlygate4sd3_1
Xhold55 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[47\] VPWR VGND
+ net98 sg13g2_dlygate4sd3_1
XFILLER_29_55 VPWR VGND sg13g2_fill_2
Xhold33 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[10\] VPWR VGND
+ net76 sg13g2_dlygate4sd3_1
Xhold44 _0134_ VPWR VGND net87 sg13g2_dlygate4sd3_1
XFILLER_48_429 VPWR VGND sg13g2_decap_8
Xhold99 _0025_ VPWR VGND net142 sg13g2_dlygate4sd3_1
Xhold66 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[66\] VPWR VGND
+ net109 sg13g2_dlygate4sd3_1
XFILLER_21_1025 VPWR VGND sg13g2_decap_4
Xhold77 _0095_ VPWR VGND net120 sg13g2_dlygate4sd3_1
Xhold88 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[13\] VPWR VGND
+ net131 sg13g2_dlygate4sd3_1
XFILLER_25_860 VPWR VGND sg13g2_fill_1
XFILLER_44_679 VPWR VGND sg13g2_decap_8
XFILLER_8_503 VPWR VGND sg13g2_fill_2
XFILLER_48_941 VPWR VGND sg13g2_decap_8
XFILLER_19_131 VPWR VGND sg13g2_decap_8
XFILLER_35_679 VPWR VGND sg13g2_fill_1
XFILLER_35_668 VPWR VGND sg13g2_decap_8
X_2952_ _1080_ VPWR _0115_ VGND net620 _1081_ sg13g2_o21ai_1
X_2883_ net834 _1034_ net740 _1037_ VPWR VGND sg13g2_nand3_1
X_4484_ net733 VGND VPWR net54 u_usb_cdc.u_sie.u_phy_rx.sample_cnt_q\[0\] clknet_leaf_30_clk_regs
+ sg13g2_dfrbpq_1
Xhold514 _1810_ VPWR VGND net557 sg13g2_dlygate4sd3_1
XFILLER_7_591 VPWR VGND sg13g2_fill_1
Xhold503 _0265_ VPWR VGND net546 sg13g2_dlygate4sd3_1
Xhold536 _0333_ VPWR VGND net855 sg13g2_dlygate4sd3_1
X_3504_ _1446_ net778 _1450_ VPWR VGND sg13g2_xor2_1
Xhold525 u_usb_cdc.u_sie.u_phy_rx.state_q\[2\] VPWR VGND net568 sg13g2_dlygate4sd3_1
X_3435_ VGND VPWR net721 net582 _0276_ _1403_ sg13g2_a21oi_1
Xhold569 u_usb_cdc.u_sie.crc16_q\[9\] VPWR VGND net888 sg13g2_dlygate4sd3_1
Xhold547 u_usb_cdc.u_ctrl_endp.req_q\[2\] VPWR VGND net866 sg13g2_dlygate4sd3_1
Xhold558 _0393_ VPWR VGND net877 sg13g2_dlygate4sd3_1
X_3366_ net755 _0601_ _1249_ _1360_ VPWR VGND sg13g2_nor3_2
X_3297_ net825 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[33\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[41\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[49\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[57\] net817 _1298_
+ VPWR VGND sg13g2_mux4_1
X_2317_ VPWR VGND _0538_ _0548_ _0536_ _0531_ _0549_ _0532_ sg13g2_a221oi_1
X_2248_ _0480_ _0479_ _0453_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_974 VPWR VGND sg13g2_decap_8
X_2179_ _1944_ net556 _2033_ VPWR VGND sg13g2_nor2_1
XFILLER_25_101 VPWR VGND sg13g2_fill_1
XFILLER_38_484 VPWR VGND sg13g2_decap_8
XFILLER_25_145 VPWR VGND sg13g2_decap_8
XFILLER_41_649 VPWR VGND sg13g2_fill_2
XFILLER_40_137 VPWR VGND sg13g2_fill_1
XFILLER_5_539 VPWR VGND sg13g2_fill_2
Xoutput23 net23 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_734 VPWR VGND sg13g2_decap_8
XFILLER_49_716 VPWR VGND sg13g2_decap_8
XFILLER_0_288 VPWR VGND sg13g2_decap_8
XFILLER_45_911 VPWR VGND sg13g2_decap_8
XFILLER_16_101 VPWR VGND sg13g2_fill_1
XFILLER_29_484 VPWR VGND sg13g2_fill_1
XFILLER_45_988 VPWR VGND sg13g2_decap_8
X_3220_ _1237_ VPWR _0227_ VGND _1915_ net603 sg13g2_o21ai_1
X_3151_ VGND VPWR _1998_ net605 _0195_ _1200_ sg13g2_a21oi_1
X_2102_ VPWR _1959_ net888 VGND sg13g2_inv_1
X_3082_ _1152_ net203 _1151_ VPWR VGND sg13g2_nand2_1
X_3984_ net748 net885 _1820_ VPWR VGND sg13g2_nor2_1
X_2935_ _1073_ VPWR _0105_ VGND net619 _1074_ sg13g2_o21ai_1
X_2866_ net4 net1006 net646 _0077_ VPWR VGND sg13g2_mux2_1
Xhold300 _1224_ VPWR VGND net343 sg13g2_dlygate4sd3_1
X_2797_ _0973_ net560 _0862_ VPWR VGND sg13g2_nand2_1
XFILLER_11_1024 VPWR VGND sg13g2_decap_4
Xhold311 u_usb_cdc.u_sie.delay_cnt_q\[0\] VPWR VGND net354 sg13g2_dlygate4sd3_1
Xhold333 u_usb_cdc.u_sie.in_byte_q\[1\] VPWR VGND net376 sg13g2_dlygate4sd3_1
Xhold322 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[1\] VPWR VGND net365 sg13g2_dlygate4sd3_1
Xhold344 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[5\] VPWR VGND net387 sg13g2_dlygate4sd3_1
Xhold366 u_usb_cdc.u_sie.addr_q\[6\] VPWR VGND net409 sg13g2_dlygate4sd3_1
Xhold355 _1177_ VPWR VGND net398 sg13g2_dlygate4sd3_1
X_4467_ net734 VGND VPWR net503 u_usb_cdc.u_sie.u_phy_rx.rx_eop_q clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_1
Xhold377 _0165_ VPWR VGND net420 sg13g2_dlygate4sd3_1
X_3418_ VGND VPWR net719 _1390_ _0267_ _1395_ sg13g2_a21oi_1
Xfanout824 net825 net824 VPWR VGND sg13g2_buf_8
Xfanout813 net1031 net813 VPWR VGND sg13g2_buf_8
Xhold399 _0184_ VPWR VGND net442 sg13g2_dlygate4sd3_1
X_4398_ net700 VGND VPWR _0326_ u_usb_cdc.u_sie.crc16_q\[3\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
Xhold388 _1479_ VPWR VGND net431 sg13g2_dlygate4sd3_1
Xfanout802 net1014 net802 VPWR VGND sg13g2_buf_8
X_3349_ _1344_ VPWR _1345_ VGND net818 net246 sg13g2_o21ai_1
Xfanout846 net1035 net846 VPWR VGND sg13g2_buf_2
Xfanout835 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] net835 VPWR VGND sg13g2_buf_8
XFILLER_45_218 VPWR VGND sg13g2_fill_2
XFILLER_27_944 VPWR VGND sg13g2_decap_8
XFILLER_45_229 VPWR VGND sg13g2_decap_4
XFILLER_42_903 VPWR VGND sg13g2_decap_8
XFILLER_26_67 VPWR VGND sg13g2_fill_2
XFILLER_13_159 VPWR VGND sg13g2_fill_1
XFILLER_1_553 VPWR VGND sg13g2_fill_2
XFILLER_49_513 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk_regs clknet_0_clk_regs clknet_3_1__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_45_752 VPWR VGND sg13g2_decap_8
XFILLER_17_498 VPWR VGND sg13g2_decap_4
XFILLER_41_991 VPWR VGND sg13g2_decap_8
X_2720_ net717 _1976_ _0916_ VPWR VGND sg13g2_nor2_1
X_2651_ _0858_ _0859_ _0860_ _0862_ VGND VPWR _0861_ sg13g2_nor4_2
XFILLER_8_196 VPWR VGND sg13g2_fill_2
X_2582_ _0805_ VPWR _0008_ VGND _0722_ _0791_ sg13g2_o21ai_1
X_4321_ net651 VGND VPWR net265 net26 clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
X_4252_ net649 VGND VPWR net223 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[14\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
X_3203_ net402 net630 _1228_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1028 VPWR VGND sg13g2_fill_1
X_4183_ net663 VGND VPWR net521 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[29\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
X_3134_ _1190_ net758 _1141_ VPWR VGND sg13g2_nand2_2
X_3065_ _1143_ net216 net634 VPWR VGND sg13g2_nand2_1
X_3967_ VGND VPWR _1944_ net708 _0399_ net533 sg13g2_a21oi_1
X_2918_ _1063_ net168 _1060_ VPWR VGND sg13g2_nand2_1
X_3898_ VGND VPWR net282 _1760_ _1766_ net879 sg13g2_a21oi_1
X_2849_ _1020_ net994 _1019_ VPWR VGND sg13g2_nand2b_1
Xhold130 _0191_ VPWR VGND net173 sg13g2_dlygate4sd3_1
Xhold152 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[27\] VPWR
+ VGND net195 sg13g2_dlygate4sd3_1
Xhold141 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[3\] VPWR VGND
+ net184 sg13g2_dlygate4sd3_1
Xhold174 _0167_ VPWR VGND net217 sg13g2_dlygate4sd3_1
Xhold163 _0119_ VPWR VGND net206 sg13g2_dlygate4sd3_1
Xhold185 u_usb_cdc.u_sie.rx_data\[4\] VPWR VGND net228 sg13g2_dlygate4sd3_1
Xfanout632 net633 net632 VPWR VGND sg13g2_buf_8
Xfanout610 net612 net610 VPWR VGND sg13g2_buf_8
Xfanout621 _1044_ net621 VPWR VGND sg13g2_buf_8
Xhold196 _0105_ VPWR VGND net239 sg13g2_dlygate4sd3_1
Xfanout676 net682 net676 VPWR VGND sg13g2_buf_8
Xfanout654 net659 net654 VPWR VGND sg13g2_buf_8
Xfanout643 _2024_ net643 VPWR VGND sg13g2_buf_8
Xfanout665 net671 net665 VPWR VGND sg13g2_buf_8
Xfanout687 net689 net687 VPWR VGND sg13g2_buf_8
Xfanout698 net699 net698 VPWR VGND sg13g2_buf_2
XFILLER_37_11 VPWR VGND sg13g2_fill_1
XFILLER_37_88 VPWR VGND sg13g2_fill_1
XFILLER_42_700 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_2_clk_regs clknet_3_1__leaf_clk_regs clknet_leaf_2_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_41_298 VPWR VGND sg13g2_decap_4
XFILLER_6_656 VPWR VGND sg13g2_decap_4
XFILLER_18_730 VPWR VGND sg13g2_fill_1
XFILLER_18_785 VPWR VGND sg13g2_fill_2
XFILLER_45_571 VPWR VGND sg13g2_fill_1
XFILLER_45_582 VPWR VGND sg13g2_fill_2
XFILLER_17_284 VPWR VGND sg13g2_fill_1
XFILLER_33_733 VPWR VGND sg13g2_decap_4
XFILLER_33_755 VPWR VGND sg13g2_fill_1
X_3821_ VGND VPWR _1709_ _1701_ _0517_ sg13g2_or2_1
X_3752_ _1653_ net866 _1568_ VPWR VGND sg13g2_nand2_1
X_2703_ _0902_ net1007 net595 VPWR VGND sg13g2_nand2b_1
X_3683_ _1586_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[67\] net628
+ VPWR VGND sg13g2_nand2_1
X_2634_ net844 net593 net750 _0845_ VPWR VGND sg13g2_nand3_1
X_2565_ _0734_ _0737_ _0717_ _0791_ VPWR VGND sg13g2_nand3_1
X_4304_ net649 VGND VPWR net208 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[66\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
X_2496_ _0723_ _0707_ _0722_ VPWR VGND sg13g2_nand2_1
X_4235_ net679 VGND VPWR net852 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[1\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
X_4166_ net662 VGND VPWR net120 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[12\]
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
X_3117_ VGND VPWR net633 _1178_ _0183_ net398 sg13g2_a21oi_1
X_4097_ net692 VGND VPWR net943 u_usb_cdc.u_ctrl_endp.req_q\[3\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_1
X_3048_ _1025_ net833 _1032_ _0160_ VPWR VGND sg13g2_mux2_1
XFILLER_36_571 VPWR VGND sg13g2_fill_1
XFILLER_12_928 VPWR VGND sg13g2_fill_2
XFILLER_11_427 VPWR VGND sg13g2_decap_4
XFILLER_11_416 VPWR VGND sg13g2_fill_2
XFILLER_2_136 VPWR VGND sg13g2_fill_1
XFILLER_24_1012 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_47_803 VPWR VGND sg13g2_decap_8
XFILLER_48_87 VPWR VGND sg13g2_fill_1
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_42_530 VPWR VGND sg13g2_decap_8
XFILLER_30_703 VPWR VGND sg13g2_fill_2
XFILLER_31_1016 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_431 VPWR VGND sg13g2_fill_2
XFILLER_7_965 VPWR VGND sg13g2_decap_8
X_2350_ _0582_ net844 _0522_ net745 net752 VPWR VGND sg13g2_a22oi_1
XFILLER_2_681 VPWR VGND sg13g2_decap_4
X_2281_ VGND VPWR _0513_ _0512_ net750 sg13g2_or2_1
X_4020_ _1851_ VPWR _1852_ VGND _2018_ _1712_ sg13g2_o21ai_1
XFILLER_29_4 VPWR VGND sg13g2_decap_8
XFILLER_49_151 VPWR VGND sg13g2_decap_4
XFILLER_49_184 VPWR VGND sg13g2_fill_2
XFILLER_18_582 VPWR VGND sg13g2_fill_2
X_3804_ _1697_ VPWR _0351_ VGND _1915_ net600 sg13g2_o21ai_1
X_3735_ _1636_ VPWR _0343_ VGND _1634_ _1635_ sg13g2_o21ai_1
X_3666_ VGND VPWR net776 _0670_ _1570_ _0647_ sg13g2_a21oi_1
X_3597_ _1503_ _1441_ net784 VPWR VGND sg13g2_nand2b_1
X_2617_ _0014_ _0832_ _0792_ VPWR VGND sg13g2_nand2b_1
XFILLER_0_629 VPWR VGND sg13g2_decap_8
XFILLER_0_607 VPWR VGND sg13g2_decap_4
X_2548_ _0775_ _0749_ _0695_ _0745_ u_usb_cdc.u_ctrl_endp.req_q\[1\] VPWR VGND sg13g2_a22oi_1
X_2479_ _0707_ u_usb_cdc.sie_out_data\[3\] _0690_ VPWR VGND sg13g2_nand2_1
X_4218_ net680 VGND VPWR net93 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[64\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
X_4149_ net661 VGND VPWR _0078_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_2
XFILLER_8_729 VPWR VGND sg13g2_decap_4
Xclkload0 clkload0/Y clknet_3_0__leaf_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_3_467 VPWR VGND sg13g2_fill_1
XFILLER_46_176 VPWR VGND sg13g2_fill_2
XFILLER_47_677 VPWR VGND sg13g2_decap_8
XFILLER_30_544 VPWR VGND sg13g2_decap_8
X_3520_ net971 net765 net587 _0306_ VPWR VGND sg13g2_mux2_1
Xhold718 u_usb_cdc.sie_in_data_ack VPWR VGND net1037 sg13g2_dlygate4sd3_1
Xhold707 u_usb_cdc.u_sie.phy_state_q\[7\] VPWR VGND net1026 sg13g2_dlygate4sd3_1
X_3451_ _1389_ _1411_ _1412_ VPWR VGND sg13g2_nor2_2
Xhold729 u_usb_cdc.rstn VPWR VGND net1048 sg13g2_dlygate4sd3_1
X_3382_ _1367_ VPWR _0258_ VGND net965 _1368_ sg13g2_o21ai_1
X_2402_ _0601_ _0617_ net968 _0632_ VPWR VGND sg13g2_nand3_1
X_2333_ _0556_ _0564_ _0565_ VPWR VGND sg13g2_nor2_1
X_2264_ _0491_ _0487_ _0496_ VPWR VGND sg13g2_xor2_1
X_2195_ _1944_ net314 net1022 _2049_ VPWR VGND _2042_ sg13g2_nand4_1
X_4003_ _1837_ _1969_ u_usb_cdc.u_sie.phy_state_q\[10\] net766 net842 VPWR VGND sg13g2_a22oi_1
XFILLER_19_891 VPWR VGND sg13g2_fill_2
XFILLER_19_880 VPWR VGND sg13g2_decap_8
XFILLER_34_850 VPWR VGND sg13g2_fill_1
XFILLER_34_883 VPWR VGND sg13g2_fill_2
X_3718_ net804 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[36\] _1620_
+ VPWR VGND sg13g2_nor2_1
X_3649_ net806 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[1\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[9\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[17\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[25\]
+ net799 _1554_ VPWR VGND sg13g2_mux4_1
XFILLER_1_905 VPWR VGND sg13g2_decap_8
Xhold23 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[10\] VPWR VGND
+ net66 sg13g2_dlygate4sd3_1
Xhold12 u_usb_cdc.u_sie.out_toggle_q\[1\] VPWR VGND net55 sg13g2_dlygate4sd3_1
Xhold56 _0214_ VPWR VGND net99 sg13g2_dlygate4sd3_1
Xhold34 _0093_ VPWR VGND net77 sg13g2_dlygate4sd3_1
Xhold45 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[48\] VPWR VGND
+ net88 sg13g2_dlygate4sd3_1
XFILLER_29_622 VPWR VGND sg13g2_fill_1
XFILLER_21_1004 VPWR VGND sg13g2_decap_8
Xhold89 _0096_ VPWR VGND net132 sg13g2_dlygate4sd3_1
Xhold67 _0149_ VPWR VGND net110 sg13g2_dlygate4sd3_1
Xhold78 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[23\] VPWR VGND
+ net121 sg13g2_dlygate4sd3_1
XFILLER_12_511 VPWR VGND sg13g2_decap_4
XFILLER_12_555 VPWR VGND sg13g2_fill_2
XFILLER_12_544 VPWR VGND sg13g2_fill_1
XFILLER_3_253 VPWR VGND sg13g2_fill_2
XFILLER_48_920 VPWR VGND sg13g2_decap_8
XFILLER_0_993 VPWR VGND sg13g2_decap_8
XFILLER_20_8 VPWR VGND sg13g2_decap_8
XFILLER_48_997 VPWR VGND sg13g2_decap_8
XFILLER_47_474 VPWR VGND sg13g2_decap_8
XFILLER_16_894 VPWR VGND sg13g2_decap_8
X_2951_ _1081_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ _1078_ VPWR VGND sg13g2_nand2_1
X_2882_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ net869 _1036_ _0090_ VPWR VGND sg13g2_mux2_1
Xhold515 _0397_ VPWR VGND net558 sg13g2_dlygate4sd3_1
X_4483_ net732 VGND VPWR net271 u_usb_cdc.u_sie.rx_data\[7\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_1
Xhold504 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q
+ VPWR VGND net547 sg13g2_dlygate4sd3_1
X_3503_ net781 net776 net785 _1449_ VPWR VGND _0540_ sg13g2_nand4_1
Xhold526 _0920_ VPWR VGND net569 sg13g2_dlygate4sd3_1
X_3434_ net485 net582 _1403_ VPWR VGND sg13g2_nor2_1
Xhold559 u_usb_cdc.addr\[5\] VPWR VGND net878 sg13g2_dlygate4sd3_1
Xhold537 u_usb_cdc.u_sie.in_toggle_q\[1\] VPWR VGND net856 sg13g2_dlygate4sd3_1
Xhold548 _0003_ VPWR VGND net867 sg13g2_dlygate4sd3_1
XFILLER_44_1026 VPWR VGND sg13g2_fill_2
X_3365_ VGND VPWR _2013_ net617 _0250_ _1359_ sg13g2_a21oi_1
X_3296_ VPWR _0243_ _1297_ VGND sg13g2_inv_1
X_2316_ net779 _0543_ _0546_ _0547_ _0548_ VPWR VGND sg13g2_nor4_1
XFILLER_39_953 VPWR VGND sg13g2_decap_8
X_2247_ _0455_ _0478_ _0479_ VPWR VGND sg13g2_and2_1
X_2178_ _2031_ VPWR _2032_ VGND u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\] _1945_ sg13g2_o21ai_1
XFILLER_26_625 VPWR VGND sg13g2_fill_2
XFILLER_5_507 VPWR VGND sg13g2_decap_8
Xoutput24 net24 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_713 VPWR VGND sg13g2_decap_8
XFILLER_0_267 VPWR VGND sg13g2_decap_8
XFILLER_48_249 VPWR VGND sg13g2_fill_2
Xclkbuf_3_0__f_clk_regs clknet_0_clk_regs clknet_3_0__leaf_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_17_614 VPWR VGND sg13g2_decap_4
XFILLER_44_422 VPWR VGND sg13g2_fill_1
XFILLER_45_967 VPWR VGND sg13g2_decap_8
XFILLER_17_669 VPWR VGND sg13g2_fill_1
XFILLER_17_658 VPWR VGND sg13g2_decap_4
XFILLER_9_813 VPWR VGND sg13g2_fill_1
XFILLER_12_396 VPWR VGND sg13g2_fill_1
XFILLER_9_846 VPWR VGND sg13g2_fill_2
XFILLER_21_90 VPWR VGND sg13g2_fill_2
XFILLER_4_595 VPWR VGND sg13g2_fill_2
X_3150_ net759 net605 _1200_ VPWR VGND sg13g2_nor2_1
XFILLER_0_790 VPWR VGND sg13g2_decap_8
X_2101_ VPWR _1958_ u_usb_cdc.u_sie.crc16_q\[10\] VGND sg13g2_inv_1
X_3081_ net831 _1140_ net739 _1151_ VPWR VGND sg13g2_nand3_1
XFILLER_39_249 VPWR VGND sg13g2_fill_2
XFILLER_48_794 VPWR VGND sg13g2_decap_8
XFILLER_23_628 VPWR VGND sg13g2_fill_1
XFILLER_22_127 VPWR VGND sg13g2_fill_1
X_3983_ _1819_ VPWR _0408_ VGND _0056_ net614 sg13g2_o21ai_1
Xclkbuf_leaf_26_clk_regs clknet_3_6__leaf_clk_regs clknet_leaf_26_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2934_ _1074_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ _1059_ VPWR VGND sg13g2_nand2_1
X_2865_ net3 net1013 net646 _0076_ VPWR VGND sg13g2_mux2_1
XFILLER_31_683 VPWR VGND sg13g2_decap_8
XFILLER_11_1003 VPWR VGND sg13g2_decap_8
Xhold301 _0216_ VPWR VGND net344 sg13g2_dlygate4sd3_1
X_2796_ VGND VPWR net55 _0971_ _0068_ _0972_ sg13g2_a21oi_1
Xhold312 _0316_ VPWR VGND net355 sg13g2_dlygate4sd3_1
Xhold334 _0320_ VPWR VGND net377 sg13g2_dlygate4sd3_1
Xhold323 _1751_ VPWR VGND net366 sg13g2_dlygate4sd3_1
Xhold367 _0312_ VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold356 _0183_ VPWR VGND net399 sg13g2_dlygate4sd3_1
X_4466_ net734 VGND VPWR _0394_ u_usb_cdc.u_sie.u_phy_rx.rx_en_q clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_2
Xhold345 _0375_ VPWR VGND net388 sg13g2_dlygate4sd3_1
Xhold378 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\] VPWR VGND net421 sg13g2_dlygate4sd3_1
X_3417_ net901 net578 _1395_ VPWR VGND sg13g2_nor2_1
Xfanout825 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[0\] net825
+ VPWR VGND sg13g2_buf_8
Xfanout814 net817 net814 VPWR VGND sg13g2_buf_8
X_4397_ net700 VGND VPWR _0325_ u_usb_cdc.u_sie.crc16_q\[2\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
Xfanout803 net806 net803 VPWR VGND sg13g2_buf_8
Xhold389 _0317_ VPWR VGND net432 sg13g2_dlygate4sd3_1
X_3348_ _1344_ net818 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[46\]
+ VPWR VGND sg13g2_nand2b_1
Xfanout836 net986 net836 VPWR VGND sg13g2_buf_8
Xfanout847 net848 net847 VPWR VGND sg13g2_buf_8
X_3279_ VGND VPWR _1278_ _1281_ _1282_ _1264_ sg13g2_a21oi_1
XFILLER_26_46 VPWR VGND sg13g2_decap_8
XFILLER_27_989 VPWR VGND sg13g2_decap_8
XFILLER_42_959 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_27_1010 VPWR VGND sg13g2_decap_8
XFILLER_49_569 VPWR VGND sg13g2_decap_8
XFILLER_37_709 VPWR VGND sg13g2_fill_2
XFILLER_44_252 VPWR VGND sg13g2_fill_2
XFILLER_33_948 VPWR VGND sg13g2_fill_1
XFILLER_41_970 VPWR VGND sg13g2_decap_8
XFILLER_9_654 VPWR VGND sg13g2_decap_4
X_2650_ _0861_ net765 u_usb_cdc.u_sie.data_q\[6\] VPWR VGND sg13g2_xnor2_1
X_2581_ net957 VPWR _0805_ VGND _0795_ _0804_ sg13g2_o21ai_1
X_4320_ net651 VGND VPWR net295 net25 clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
XFILLER_5_882 VPWR VGND sg13g2_decap_4
X_4251_ net658 VGND VPWR net269 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[13\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_3202_ VGND VPWR _1915_ net630 _0219_ _1227_ sg13g2_a21oi_1
X_4182_ net663 VGND VPWR net536 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[28\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
X_3133_ net345 net632 _1189_ VPWR VGND sg13g2_nor2_1
X_3064_ _1140_ net739 _1142_ VPWR VGND net831 sg13g2_nand3b_1
XFILLER_48_591 VPWR VGND sg13g2_decap_8
X_3966_ net532 net708 _1812_ VPWR VGND sg13g2_nor2_1
X_2917_ _1061_ VPWR _0099_ VGND net620 _1062_ sg13g2_o21ai_1
XFILLER_31_491 VPWR VGND sg13g2_decap_8
X_3897_ _1765_ net282 net879 _1760_ VPWR VGND sg13g2_and3_1
X_2848_ net834 net833 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\]
+ _1019_ VPWR VGND sg13g2_nor3_2
X_2779_ net768 _0952_ _0956_ _0957_ VPWR VGND sg13g2_nor3_1
Xhold120 _0212_ VPWR VGND net163 sg13g2_dlygate4sd3_1
Xhold142 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[36\] VPWR
+ VGND net185 sg13g2_dlygate4sd3_1
Xhold153 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[38\] VPWR VGND
+ net196 sg13g2_dlygate4sd3_1
Xhold131 _0052_ VPWR VGND net174 sg13g2_dlygate4sd3_1
Xhold164 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[66\] VPWR
+ VGND net207 sg13g2_dlygate4sd3_1
Xhold186 _0405_ VPWR VGND net229 sg13g2_dlygate4sd3_1
Xhold175 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[33\] VPWR VGND
+ net218 sg13g2_dlygate4sd3_1
X_4449_ net725 VGND VPWR _0377_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[7\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
Xfanout633 _1176_ net633 VPWR VGND sg13g2_buf_8
Xfanout600 net602 net600 VPWR VGND sg13g2_buf_8
Xfanout622 net623 net622 VPWR VGND sg13g2_buf_8
Xfanout611 net612 net611 VPWR VGND sg13g2_buf_2
Xhold197 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[53\] VPWR VGND
+ net240 sg13g2_dlygate4sd3_1
Xfanout655 net659 net655 VPWR VGND sg13g2_buf_8
Xfanout666 net667 net666 VPWR VGND sg13g2_buf_8
Xfanout644 _1059_ net644 VPWR VGND sg13g2_buf_8
Xfanout677 net682 net677 VPWR VGND sg13g2_buf_8
Xfanout688 net689 net688 VPWR VGND sg13g2_buf_1
Xfanout699 net704 net699 VPWR VGND sg13g2_buf_8
XFILLER_37_67 VPWR VGND sg13g2_decap_4
XFILLER_46_539 VPWR VGND sg13g2_fill_1
XFILLER_27_742 VPWR VGND sg13g2_decap_8
XFILLER_15_915 VPWR VGND sg13g2_fill_2
XFILLER_41_233 VPWR VGND sg13g2_fill_2
XFILLER_30_907 VPWR VGND sg13g2_fill_1
XFILLER_23_992 VPWR VGND sg13g2_decap_8
XFILLER_10_642 VPWR VGND sg13g2_fill_2
XFILLER_1_395 VPWR VGND sg13g2_decap_8
XFILLER_49_344 VPWR VGND sg13g2_decap_8
XFILLER_18_764 VPWR VGND sg13g2_fill_1
X_3820_ _1708_ net944 _1703_ _0356_ VPWR VGND sg13g2_mux2_1
X_3751_ _1926_ _0533_ _0657_ _1652_ VPWR VGND sg13g2_or3_1
X_2702_ VGND VPWR net707 _0901_ _0900_ net976 sg13g2_a21oi_2
X_3682_ _1585_ VPWR _0341_ VGND _1583_ _1584_ sg13g2_o21ai_1
X_2633_ _0844_ net750 net593 VPWR VGND sg13g2_nand2_1
X_2564_ net513 VPWR _0790_ VGND _0704_ _0789_ sg13g2_o21ai_1
X_4303_ net650 VGND VPWR net130 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[65\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
X_2495_ u_usb_cdc.sie_out_data\[2\] _0689_ net720 _0722_ VPWR VGND sg13g2_nand3_1
X_4234_ net681 VGND VPWR _0163_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[0\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_2
X_4165_ net660 VGND VPWR net79 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[11\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
X_3116_ _1178_ net764 _1141_ VPWR VGND sg13g2_nand2_2
Xclkbuf_leaf_41_clk_regs clknet_3_5__leaf_clk_regs clknet_leaf_41_clk_regs VPWR VGND
+ sg13g2_buf_8
X_4096_ net693 VGND VPWR net867 u_usb_cdc.u_ctrl_endp.req_q\[2\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
X_3047_ _1023_ net977 _1032_ _0159_ VPWR VGND sg13g2_mux2_1
XFILLER_36_594 VPWR VGND sg13g2_fill_2
XFILLER_17_1020 VPWR VGND sg13g2_decap_8
X_3949_ VGND VPWR net744 net387 _1803_ net917 sg13g2_a21oi_1
XFILLER_20_973 VPWR VGND sg13g2_fill_2
XFILLER_47_859 VPWR VGND sg13g2_decap_8
XFILLER_15_734 VPWR VGND sg13g2_fill_2
XFILLER_30_737 VPWR VGND sg13g2_decap_4
XFILLER_6_465 VPWR VGND sg13g2_decap_4
XFILLER_6_498 VPWR VGND sg13g2_decap_4
XFILLER_2_660 VPWR VGND sg13g2_decap_8
X_2280_ _0512_ net841 _0510_ VPWR VGND sg13g2_nand2_1
XFILLER_38_804 VPWR VGND sg13g2_fill_1
XFILLER_49_196 VPWR VGND sg13g2_decap_8
X_3803_ net592 _1692_ net997 _1697_ VPWR VGND sg13g2_nand3_1
XFILLER_20_258 VPWR VGND sg13g2_fill_1
X_3734_ _1636_ net997 net597 VPWR VGND sg13g2_nand2_1
X_3665_ net773 _1568_ _1569_ VPWR VGND sg13g2_nor2_1
X_2616_ _0832_ _0827_ net1030 _0822_ _0667_ VPWR VGND sg13g2_a22oi_1
XFILLER_47_1013 VPWR VGND sg13g2_decap_8
X_3596_ _0652_ _1501_ _1502_ VPWR VGND sg13g2_nor2_1
X_2547_ _0672_ _0773_ _0774_ VPWR VGND sg13g2_nor2_1
X_2478_ _0706_ u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] VPWR VGND net413 sg13g2_nand2b_2
X_4217_ net669 VGND VPWR net478 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[63\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_4148_ net661 VGND VPWR _0077_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_2
XFILLER_37_870 VPWR VGND sg13g2_fill_1
X_4079_ net598 _0586_ _1524_ _1899_ VPWR VGND sg13g2_nor3_1
XFILLER_24_542 VPWR VGND sg13g2_fill_2
XFILLER_11_236 VPWR VGND sg13g2_fill_2
Xclkload1 clknet_3_7__leaf_clk_regs clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_47_656 VPWR VGND sg13g2_decap_8
XFILLER_43_884 VPWR VGND sg13g2_decap_8
XFILLER_15_586 VPWR VGND sg13g2_fill_1
XFILLER_30_501 VPWR VGND sg13g2_fill_2
XFILLER_7_730 VPWR VGND sg13g2_fill_1
XFILLER_11_792 VPWR VGND sg13g2_fill_1
Xhold708 _0875_ VPWR VGND net1027 sg13g2_dlygate4sd3_1
Xhold719 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[0\] VPWR VGND
+ net1038 sg13g2_dlygate4sd3_1
X_3450_ VGND VPWR _0634_ _0685_ _1411_ net624 sg13g2_a21oi_1
X_3381_ VGND VPWR _1368_ _1365_ net617 sg13g2_or2_1
X_2401_ _0611_ _0616_ net624 _0631_ VPWR VGND sg13g2_nor3_1
X_2332_ net710 VPWR _0564_ VGND _0561_ _0563_ sg13g2_o21ai_1
X_2263_ _0494_ _0491_ _0495_ VPWR VGND sg13g2_xor2_1
X_4002_ net625 VPWR _1836_ VGND net439 _1835_ sg13g2_o21ai_1
X_2194_ _2039_ _2042_ net961 _2048_ VPWR VGND _2047_ sg13g2_nand4_1
XFILLER_26_818 VPWR VGND sg13g2_fill_1
XFILLER_37_177 VPWR VGND sg13g2_fill_1
XFILLER_21_578 VPWR VGND sg13g2_decap_4
X_3717_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[44\] net805 _1619_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_20_15 VPWR VGND sg13g2_decap_4
X_3648_ _1553_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[65\] net628
+ VPWR VGND sg13g2_nand2_1
X_3579_ _0328_ net579 _0489_ net583 _1966_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_449 VPWR VGND sg13g2_decap_8
Xhold13 _0068_ VPWR VGND net56 sg13g2_dlygate4sd3_1
XFILLER_48_409 VPWR VGND sg13g2_decap_4
Xhold24 _0177_ VPWR VGND net67 sg13g2_dlygate4sd3_1
Xhold35 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[11\] VPWR VGND
+ net78 sg13g2_dlygate4sd3_1
Xhold46 _0131_ VPWR VGND net89 sg13g2_dlygate4sd3_1
XFILLER_29_601 VPWR VGND sg13g2_decap_8
Xhold57 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[57\] VPWR VGND
+ net100 sg13g2_dlygate4sd3_1
Xhold68 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[12\] VPWR VGND
+ net111 sg13g2_dlygate4sd3_1
Xhold79 _0106_ VPWR VGND net122 sg13g2_dlygate4sd3_1
XFILLER_12_567 VPWR VGND sg13g2_fill_1
XFILLER_12_578 VPWR VGND sg13g2_decap_8
XFILLER_4_711 VPWR VGND sg13g2_fill_2
XFILLER_0_972 VPWR VGND sg13g2_decap_8
XFILLER_39_409 VPWR VGND sg13g2_decap_8
XFILLER_48_976 VPWR VGND sg13g2_decap_8
XFILLER_47_464 VPWR VGND sg13g2_decap_4
XFILLER_35_648 VPWR VGND sg13g2_decap_8
X_2950_ _1080_ net158 _1079_ VPWR VGND sg13g2_nand2_1
X_2881_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net526 _1036_ _0089_ VPWR VGND sg13g2_mux2_1
XFILLER_42_180 VPWR VGND sg13g2_fill_2
XFILLER_7_582 VPWR VGND sg13g2_fill_2
Xhold516 u_usb_cdc.u_ctrl_endp.addr_dd\[3\] VPWR VGND net559 sg13g2_dlygate4sd3_1
X_4482_ net730 VGND VPWR _0407_ u_usb_cdc.u_sie.rx_data\[6\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_1
Xhold527 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[30\] VPWR VGND
+ net570 sg13g2_dlygate4sd3_1
Xhold505 _0074_ VPWR VGND net548 sg13g2_dlygate4sd3_1
X_3502_ _1448_ net778 _1437_ VPWR VGND sg13g2_nand2_1
Xhold549 u_usb_cdc.addr\[0\] VPWR VGND net868 sg13g2_dlygate4sd3_1
X_3433_ VGND VPWR net724 net582 _0275_ _1402_ sg13g2_a21oi_1
Xhold538 _0993_ VPWR VGND net857 sg13g2_dlygate4sd3_1
XFILLER_44_1005 VPWR VGND sg13g2_decap_8
X_3364_ VPWR VGND _1983_ net617 _1358_ net170 _1359_ _1294_ sg13g2_a221oi_1
X_3295_ _1296_ VPWR _1297_ VGND net985 _1283_ sg13g2_o21ai_1
X_2315_ _0547_ net772 u_usb_cdc.u_ctrl_endp.req_q\[8\] VPWR VGND sg13g2_nand2_1
X_2246_ _0463_ _0473_ _0474_ _0477_ _0478_ VPWR VGND sg13g2_and4_1
X_2177_ _2031_ _1943_ net553 VPWR VGND sg13g2_nand2_1
XFILLER_31_58 VPWR VGND sg13g2_decap_8
Xoutput25 net25 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput14 net14 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_769 VPWR VGND sg13g2_decap_8
XFILLER_0_246 VPWR VGND sg13g2_decap_8
XFILLER_45_946 VPWR VGND sg13g2_decap_8
XFILLER_12_342 VPWR VGND sg13g2_decap_8
XFILLER_12_353 VPWR VGND sg13g2_fill_1
XFILLER_9_836 VPWR VGND sg13g2_fill_1
XFILLER_8_368 VPWR VGND sg13g2_fill_1
XFILLER_4_530 VPWR VGND sg13g2_fill_1
X_2100_ VPWR _1957_ u_usb_cdc.u_sie.crc16_q\[11\] VGND sg13g2_inv_1
X_3080_ _1150_ VPWR _0174_ VGND net719 net635 sg13g2_o21ai_1
XFILLER_36_902 VPWR VGND sg13g2_fill_2
XFILLER_48_773 VPWR VGND sg13g2_decap_8
XFILLER_23_618 VPWR VGND sg13g2_fill_2
X_3982_ _1819_ net270 net614 VPWR VGND sg13g2_nand2_1
XFILLER_16_692 VPWR VGND sg13g2_fill_2
X_2933_ _1073_ net238 _1060_ VPWR VGND sg13g2_nand2_1
X_2864_ net2 net1018 net646 _0075_ VPWR VGND sg13g2_mux2_1
X_2795_ _0965_ VPWR _0972_ VGND net55 _0971_ sg13g2_o21ai_1
Xhold302 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[22\] VPWR
+ VGND net345 sg13g2_dlygate4sd3_1
Xhold335 u_usb_cdc.u_sie.in_toggle_q\[2\] VPWR VGND net378 sg13g2_dlygate4sd3_1
Xhold313 u_usb_cdc.u_sie.u_phy_tx.data_q\[5\] VPWR VGND net356 sg13g2_dlygate4sd3_1
Xhold324 _0371_ VPWR VGND net367 sg13g2_dlygate4sd3_1
Xhold368 u_usb_cdc.u_ctrl_endp.req_q\[10\] VPWR VGND net411 sg13g2_dlygate4sd3_1
Xhold357 u_usb_cdc.u_sie.in_byte_q\[3\] VPWR VGND net400 sg13g2_dlygate4sd3_1
X_4465_ net734 VGND VPWR net877 u_usb_cdc.u_sie.rx_err clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
Xhold346 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[1\] VPWR VGND net389 sg13g2_dlygate4sd3_1
Xhold379 _0363_ VPWR VGND net422 sg13g2_dlygate4sd3_1
X_3416_ VGND VPWR net720 net578 _0266_ _1394_ sg13g2_a21oi_1
Xfanout815 net817 net815 VPWR VGND sg13g2_buf_1
X_4396_ net695 VGND VPWR _0324_ u_usb_cdc.u_sie.crc16_q\[1\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xfanout804 net806 net804 VPWR VGND sg13g2_buf_8
Xfanout826 net1042 net826 VPWR VGND sg13g2_buf_8
X_3347_ VGND VPWR net815 _1342_ _1343_ net813 sg13g2_a21oi_1
Xfanout848 net1047 net848 VPWR VGND sg13g2_buf_2
Xfanout837 u_usb_cdc.u_sie.phy_state_q\[10\] net837 VPWR VGND sg13g2_buf_8
X_3278_ _1281_ _0604_ _1280_ net951 net755 VPWR VGND sg13g2_a22oi_1
XFILLER_27_902 VPWR VGND sg13g2_decap_4
X_2229_ _0461_ _0459_ _0460_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_27_968 VPWR VGND sg13g2_decap_8
XFILLER_42_938 VPWR VGND sg13g2_decap_8
XFILLER_26_69 VPWR VGND sg13g2_fill_1
XFILLER_35_990 VPWR VGND sg13g2_decap_8
XFILLER_13_128 VPWR VGND sg13g2_fill_2
XFILLER_22_651 VPWR VGND sg13g2_decap_4
XFILLER_42_35 VPWR VGND sg13g2_fill_2
XFILLER_22_695 VPWR VGND sg13g2_fill_2
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_4
XFILLER_49_548 VPWR VGND sg13g2_decap_8
XFILLER_18_924 VPWR VGND sg13g2_fill_1
XFILLER_29_283 VPWR VGND sg13g2_fill_2
XFILLER_45_787 VPWR VGND sg13g2_decap_8
XFILLER_34_1015 VPWR VGND sg13g2_decap_8
X_2580_ _0796_ _0803_ _0699_ _0804_ VPWR VGND sg13g2_nand3_1
XFILLER_8_198 VPWR VGND sg13g2_fill_1
X_4250_ net654 VGND VPWR net112 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[12\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_3201_ net498 net630 _1227_ VPWR VGND sg13g2_nor2_1
X_4181_ net665 VGND VPWR net529 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[27\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
XFILLER_41_1019 VPWR VGND sg13g2_decap_8
X_3132_ VGND VPWR net633 _1188_ _0188_ net359 sg13g2_a21oi_1
X_3063_ _1141_ net711 _1139_ VPWR VGND sg13g2_nand2_2
X_3965_ VGND VPWR _1943_ net708 _0398_ net453 sg13g2_a21oi_1
X_2916_ _1062_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net644 VPWR VGND sg13g2_nand2_1
XFILLER_32_982 VPWR VGND sg13g2_decap_8
X_3896_ VGND VPWR net282 _1762_ _0376_ _1764_ sg13g2_a21oi_1
X_2847_ net834 net833 _1018_ VPWR VGND sg13g2_nor2_1
Xhold110 _0231_ VPWR VGND net153 sg13g2_dlygate4sd3_1
X_2778_ _0956_ net710 _0955_ VPWR VGND sg13g2_nand2_2
Xhold132 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[42\] VPWR
+ VGND net175 sg13g2_dlygate4sd3_1
Xhold143 _0203_ VPWR VGND net186 sg13g2_dlygate4sd3_1
Xhold121 u_usb_cdc.u_sie.in_zlp_q\[0\] VPWR VGND net164 sg13g2_dlygate4sd3_1
Xhold165 _0233_ VPWR VGND net208 sg13g2_dlygate4sd3_1
Xhold176 _0116_ VPWR VGND net219 sg13g2_dlygate4sd3_1
Xhold154 _0121_ VPWR VGND net197 sg13g2_dlygate4sd3_1
X_4448_ net725 VGND VPWR net283 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[6\] clknet_leaf_23_clk_regs
+ sg13g2_dfrbpq_1
Xfanout623 _0697_ net623 VPWR VGND sg13g2_buf_8
Xhold187 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[44\] VPWR
+ VGND net230 sg13g2_dlygate4sd3_1
Xfanout601 net602 net601 VPWR VGND sg13g2_buf_1
Xhold198 _0136_ VPWR VGND net241 sg13g2_dlygate4sd3_1
Xfanout612 _1099_ net612 VPWR VGND sg13g2_buf_8
X_4379_ net677 VGND VPWR _0307_ u_usb_cdc.u_sie.addr_q\[1\] clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_1
Xfanout656 net659 net656 VPWR VGND sg13g2_buf_8
Xfanout634 net635 net634 VPWR VGND sg13g2_buf_8
Xfanout667 net671 net667 VPWR VGND sg13g2_buf_8
Xfanout645 _1039_ net645 VPWR VGND sg13g2_buf_8
Xfanout689 net690 net689 VPWR VGND sg13g2_buf_8
Xfanout678 net680 net678 VPWR VGND sg13g2_buf_8
XFILLER_2_1024 VPWR VGND sg13g2_decap_4
XFILLER_15_905 VPWR VGND sg13g2_decap_4
XFILLER_27_776 VPWR VGND sg13g2_fill_2
XFILLER_27_787 VPWR VGND sg13g2_fill_1
XFILLER_27_798 VPWR VGND sg13g2_fill_1
XFILLER_30_919 VPWR VGND sg13g2_decap_8
XFILLER_1_374 VPWR VGND sg13g2_decap_8
XFILLER_49_367 VPWR VGND sg13g2_fill_2
XFILLER_49_378 VPWR VGND sg13g2_decap_8
XFILLER_45_584 VPWR VGND sg13g2_fill_1
X_3750_ _1638_ VPWR _1651_ VGND net795 _1650_ sg13g2_o21ai_1
X_2701_ VPWR _0900_ _0899_ VGND sg13g2_inv_1
X_3681_ _1585_ net519 net597 VPWR VGND sg13g2_nand2_1
X_2632_ _0843_ net524 net596 VPWR VGND sg13g2_nand2_1
X_2563_ _0786_ _0788_ _0680_ _0789_ VPWR VGND sg13g2_nand3_1
X_4302_ net648 VGND VPWR net153 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[64\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
X_2494_ _0721_ net942 _0679_ VPWR VGND sg13g2_nand2_1
X_4233_ net679 VGND VPWR _0162_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_2
X_4164_ net660 VGND VPWR net77 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[10\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_1
X_4095_ net686 VGND VPWR net895 u_usb_cdc.u_ctrl_endp.req_q\[1\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_2
X_3115_ net397 net633 _1177_ VPWR VGND sg13g2_nor2_1
X_3046_ VPWR _0158_ _1132_ VGND sg13g2_inv_1
XFILLER_24_746 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_10_clk_regs clknet_3_2__leaf_clk_regs clknet_leaf_10_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3948_ net713 _1744_ _1802_ VPWR VGND sg13g2_nor2_1
X_3879_ net336 VPWR _1752_ VGND net716 _1749_ sg13g2_o21ai_1
XFILLER_3_606 VPWR VGND sg13g2_fill_1
XFILLER_48_56 VPWR VGND sg13g2_fill_2
XFILLER_47_838 VPWR VGND sg13g2_decap_8
XFILLER_48_78 VPWR VGND sg13g2_decap_8
XFILLER_15_757 VPWR VGND sg13g2_decap_4
XFILLER_6_433 VPWR VGND sg13g2_fill_1
XFILLER_11_996 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_fill_1
XFILLER_21_705 VPWR VGND sg13g2_decap_8
X_3802_ _1696_ VPWR _0350_ VGND _1912_ net600 sg13g2_o21ai_1
X_3733_ net602 VPWR _1635_ VGND net228 _1523_ sg13g2_o21ai_1
X_3664_ net792 _0533_ _0657_ _1568_ VPWR VGND sg13g2_nor3_1
X_2615_ _0013_ _0830_ _0831_ VPWR VGND sg13g2_nand2_1
X_3595_ VGND VPWR net784 _0675_ _1501_ net783 sg13g2_a21oi_1
X_2546_ VPWR VGND u_usb_cdc.u_ctrl_endp.req_q\[1\] _0772_ _0771_ u_usb_cdc.u_ctrl_endp.req_q\[11\]
+ _0773_ _0693_ sg13g2_a221oi_1
X_2477_ net874 VPWR _0705_ VGND _0696_ _0704_ sg13g2_o21ai_1
X_4216_ net668 VGND VPWR net480 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[62\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_4147_ net661 VGND VPWR _0076_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_2
X_4078_ _1896_ VPWR _0424_ VGND _1892_ _1898_ sg13g2_o21ai_1
X_3029_ _1123_ net133 _1118_ VPWR VGND sg13g2_nand2_1
Xclkload2 VPWR clkload2/Y clknet_leaf_38_clk_regs VGND sg13g2_inv_1
XFILLER_47_613 VPWR VGND sg13g2_fill_1
XFILLER_47_635 VPWR VGND sg13g2_decap_8
XFILLER_15_576 VPWR VGND sg13g2_fill_2
Xhold709 u_usb_cdc.u_sie.pid_q\[3\] VPWR VGND net1028 sg13g2_dlygate4sd3_1
X_2400_ _0630_ net850 _0601_ VPWR VGND sg13g2_nand2_2
X_3380_ net965 VPWR _1367_ VGND net617 _1366_ sg13g2_o21ai_1
X_2331_ _0559_ _0562_ _0557_ _0563_ VPWR VGND sg13g2_nand3_1
X_2262_ _0494_ _0492_ _0493_ VPWR VGND sg13g2_xnor2_1
X_4001_ _2027_ _1008_ _1835_ VPWR VGND sg13g2_nor2_1
X_2193_ _1943_ _2045_ _0056_ _2047_ VPWR VGND _2046_ sg13g2_nand4_1
XFILLER_38_635 VPWR VGND sg13g2_decap_4
XFILLER_38_679 VPWR VGND sg13g2_fill_2
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_46_690 VPWR VGND sg13g2_decap_8
XFILLER_21_513 VPWR VGND sg13g2_fill_1
X_3716_ _1617_ VPWR _1618_ VGND net798 _1615_ sg13g2_o21ai_1
X_3647_ _1549_ VPWR _1552_ VGND _1550_ _1551_ sg13g2_o21ai_1
X_3578_ _0327_ net579 _0505_ net583 _1967_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_428 VPWR VGND sg13g2_decap_8
X_2529_ _0746_ _0755_ _0743_ _0756_ VPWR VGND sg13g2_nand3_1
Xhold14 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[2\] VPWR VGND net57 sg13g2_dlygate4sd3_1
XFILLER_29_25 VPWR VGND sg13g2_decap_8
Xhold36 _0094_ VPWR VGND net79 sg13g2_dlygate4sd3_1
Xhold47 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[44\] VPWR VGND
+ net90 sg13g2_dlygate4sd3_1
Xhold25 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[70\] VPWR VGND
+ net68 sg13g2_dlygate4sd3_1
Xhold58 _1234_ VPWR VGND net101 sg13g2_dlygate4sd3_1
Xhold69 _0179_ VPWR VGND net112 sg13g2_dlygate4sd3_1
XFILLER_29_635 VPWR VGND sg13g2_decap_8
XFILLER_28_167 VPWR VGND sg13g2_decap_4
XFILLER_25_874 VPWR VGND sg13g2_fill_1
XFILLER_12_524 VPWR VGND sg13g2_fill_2
XFILLER_12_557 VPWR VGND sg13g2_fill_1
XFILLER_3_233 VPWR VGND sg13g2_fill_2
XFILLER_4_767 VPWR VGND sg13g2_fill_2
XFILLER_3_255 VPWR VGND sg13g2_fill_1
XFILLER_0_951 VPWR VGND sg13g2_decap_8
XFILLER_48_955 VPWR VGND sg13g2_decap_8
XFILLER_47_432 VPWR VGND sg13g2_fill_2
XFILLER_19_156 VPWR VGND sg13g2_fill_2
XFILLER_47_443 VPWR VGND sg13g2_decap_8
XFILLER_37_1013 VPWR VGND sg13g2_decap_8
X_2880_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net455 _1036_ _0088_ VPWR VGND sg13g2_mux2_1
XFILLER_43_682 VPWR VGND sg13g2_fill_1
Xhold506 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[1\] VPWR VGND
+ net549 sg13g2_dlygate4sd3_1
Xhold517 u_usb_cdc.u_sie.data_q\[1\] VPWR VGND net560 sg13g2_dlygate4sd3_1
X_4481_ net729 VGND VPWR net237 u_usb_cdc.u_sie.rx_data\[5\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_1
X_3501_ _1445_ VPWR _0298_ VGND _1439_ _1447_ sg13g2_o21ai_1
X_3432_ net499 net582 _1402_ VPWR VGND sg13g2_nor2_1
Xhold539 _0070_ VPWR VGND net858 sg13g2_dlygate4sd3_1
Xhold528 _0113_ VPWR VGND net571 sg13g2_dlygate4sd3_1
X_3363_ _1357_ VPWR _1358_ VGND _1288_ _1354_ sg13g2_o21ai_1
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
X_3294_ _1295_ VPWR _1296_ VGND net965 _1293_ sg13g2_o21ai_1
X_2314_ VGND VPWR _0546_ net775 net776 sg13g2_or2_1
X_2245_ _0476_ VPWR _0477_ VGND u_usb_cdc.u_sie.data_q\[6\] _0475_ sg13g2_o21ai_1
XFILLER_39_988 VPWR VGND sg13g2_decap_8
X_2176_ _0065_ net717 _2006_ VPWR VGND sg13g2_nand2_1
XFILLER_38_498 VPWR VGND sg13g2_fill_2
XFILLER_25_137 VPWR VGND sg13g2_fill_2
XFILLER_25_159 VPWR VGND sg13g2_fill_1
XFILLER_41_619 VPWR VGND sg13g2_decap_4
XFILLER_22_899 VPWR VGND sg13g2_fill_2
Xoutput15 net15 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput26 net26 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_748 VPWR VGND sg13g2_decap_8
XFILLER_0_225 VPWR VGND sg13g2_decap_8
XFILLER_45_925 VPWR VGND sg13g2_decap_8
XFILLER_17_627 VPWR VGND sg13g2_decap_4
XFILLER_8_347 VPWR VGND sg13g2_fill_2
XFILLER_21_92 VPWR VGND sg13g2_fill_1
XFILLER_4_597 VPWR VGND sg13g2_fill_1
XFILLER_47_240 VPWR VGND sg13g2_fill_2
XFILLER_48_752 VPWR VGND sg13g2_decap_8
X_3981_ net496 net506 net614 _0407_ VPWR VGND sg13g2_mux2_1
XFILLER_44_991 VPWR VGND sg13g2_decap_8
X_2932_ _1071_ VPWR _0104_ VGND net619 _1072_ sg13g2_o21ai_1
XFILLER_31_652 VPWR VGND sg13g2_fill_2
X_2863_ _0074_ net647 _1033_ VPWR VGND sg13g2_nand2_1
X_2794_ _0966_ _0969_ _0970_ _0971_ VPWR VGND sg13g2_nor3_1
Xhold303 _0189_ VPWR VGND net346 sg13g2_dlygate4sd3_1
Xhold314 _0415_ VPWR VGND net357 sg13g2_dlygate4sd3_1
Xhold325 _0053_ VPWR VGND net368 sg13g2_dlygate4sd3_1
Xhold336 _0998_ VPWR VGND net379 sg13g2_dlygate4sd3_1
Xhold369 _0000_ VPWR VGND net412 sg13g2_dlygate4sd3_1
Xhold347 _0423_ VPWR VGND net390 sg13g2_dlygate4sd3_1
Xhold358 _0322_ VPWR VGND net401 sg13g2_dlygate4sd3_1
X_4464_ net734 VGND VPWR net466 u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_1
X_3415_ net500 net578 _1394_ VPWR VGND sg13g2_nor2_1
Xfanout816 net817 net816 VPWR VGND sg13g2_buf_8
X_4395_ net695 VGND VPWR net531 u_usb_cdc.u_sie.crc16_q\[0\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_35_clk_regs clknet_3_5__leaf_clk_regs clknet_leaf_35_clk_regs VPWR VGND
+ sg13g2_buf_8
Xfanout805 net806 net805 VPWR VGND sg13g2_buf_1
X_3346_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[22\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[30\]
+ net818 _1342_ VPWR VGND sg13g2_mux2_1
Xfanout827 net828 net827 VPWR VGND sg13g2_buf_8
Xfanout838 u_usb_cdc.u_sie.phy_state_q\[9\] net838 VPWR VGND sg13g2_buf_8
Xfanout849 net969 net849 VPWR VGND sg13g2_buf_8
X_3277_ _1279_ VPWR _1280_ VGND net770 _1981_ sg13g2_o21ai_1
X_2228_ _0460_ net760 net758 VPWR VGND sg13g2_xnor2_1
X_2159_ net995 net971 net972 _2015_ VPWR VGND sg13g2_nor3_2
XFILLER_42_917 VPWR VGND sg13g2_decap_8
XFILLER_41_405 VPWR VGND sg13g2_decap_4
XFILLER_22_630 VPWR VGND sg13g2_decap_8
XFILLER_49_527 VPWR VGND sg13g2_decap_8
XFILLER_18_958 VPWR VGND sg13g2_decap_4
XFILLER_44_254 VPWR VGND sg13g2_fill_1
XFILLER_45_766 VPWR VGND sg13g2_decap_8
XFILLER_4_383 VPWR VGND sg13g2_fill_2
X_3200_ VGND VPWR net720 net630 _0218_ _1226_ sg13g2_a21oi_1
X_4180_ net660 VGND VPWR net538 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[26\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_1
X_3131_ _1188_ u_usb_cdc.sie_out_data\[5\] _1141_ VPWR VGND sg13g2_nand2_2
X_3062_ net829 net827 net826 _1140_ VPWR VGND sg13g2_nor3_1
XFILLER_36_733 VPWR VGND sg13g2_fill_2
X_3964_ net452 net708 _1811_ VPWR VGND sg13g2_nor2_1
X_2915_ _1061_ net250 _1060_ VPWR VGND sg13g2_nand2_1
X_3895_ VGND VPWR net615 _1760_ _1764_ net282 sg13g2_a21oi_1
X_2846_ _1985_ _1016_ _1017_ VPWR VGND sg13g2_nor2_1
Xhold100 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[33\] VPWR
+ VGND net143 sg13g2_dlygate4sd3_1
X_2777_ _0955_ u_usb_cdc.u_sie.pid_q\[3\] _0954_ VPWR VGND sg13g2_xnor2_1
Xhold133 _0209_ VPWR VGND net176 sg13g2_dlygate4sd3_1
Xhold111 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[34\] VPWR VGND
+ net154 sg13g2_dlygate4sd3_1
Xhold144 u_usb_cdc.u_sie.rx_data\[0\] VPWR VGND net187 sg13g2_dlygate4sd3_1
Xhold122 _0426_ VPWR VGND net165 sg13g2_dlygate4sd3_1
X_4516_ net679 VGND VPWR _0428_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
Xhold166 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[2\] VPWR VGND net209 sg13g2_dlygate4sd3_1
Xhold177 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[14\] VPWR VGND
+ net220 sg13g2_dlygate4sd3_1
Xhold155 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[35\] VPWR VGND
+ net198 sg13g2_dlygate4sd3_1
X_4447_ net725 VGND VPWR net388 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[5\] clknet_leaf_23_clk_regs
+ sg13g2_dfrbpq_1
Xhold188 _0211_ VPWR VGND net231 sg13g2_dlygate4sd3_1
Xfanout624 _0630_ net624 VPWR VGND sg13g2_buf_8
Xfanout602 _0439_ net602 VPWR VGND sg13g2_buf_8
Xfanout613 net614 net613 VPWR VGND sg13g2_buf_8
Xhold199 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[54\] VPWR VGND
+ net242 sg13g2_dlygate4sd3_1
X_4378_ net688 VGND VPWR _0306_ u_usb_cdc.endp\[3\] clknet_leaf_42_clk_regs sg13g2_dfrbpq_2
Xfanout635 _1142_ net635 VPWR VGND sg13g2_buf_8
Xfanout657 net659 net657 VPWR VGND sg13g2_buf_8
Xfanout646 net647 net646 VPWR VGND sg13g2_buf_8
X_3329_ VGND VPWR _1327_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[20\]
+ net823 sg13g2_or2_1
Xfanout668 net670 net668 VPWR VGND sg13g2_buf_8
Xfanout679 net680 net679 VPWR VGND sg13g2_buf_8
XFILLER_2_1003 VPWR VGND sg13g2_decap_8
XFILLER_41_235 VPWR VGND sg13g2_fill_1
XFILLER_6_626 VPWR VGND sg13g2_decap_8
XFILLER_1_353 VPWR VGND sg13g2_decap_8
XFILLER_40_1020 VPWR VGND sg13g2_decap_4
XFILLER_18_744 VPWR VGND sg13g2_fill_1
XFILLER_33_769 VPWR VGND sg13g2_fill_2
XFILLER_21_909 VPWR VGND sg13g2_fill_1
X_2700_ _2032_ _2037_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] _0899_ VPWR VGND _0898_
+ sg13g2_nand4_1
X_3680_ net602 VPWR _1584_ VGND net232 _1523_ sg13g2_o21ai_1
X_2631_ _0840_ VPWR _0020_ VGND _0841_ _0842_ sg13g2_o21ai_1
X_2562_ _0788_ _0631_ _0787_ VPWR VGND sg13g2_nand2_1
X_4301_ net658 VGND VPWR net149 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[63\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_2493_ _0705_ VPWR _0005_ VGND _0711_ _0720_ sg13g2_o21ai_1
X_4232_ net679 VGND VPWR _0161_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_2
X_4163_ net660 VGND VPWR net194 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[9\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_1
X_3114_ net827 net1054 _1175_ _1176_ VPWR VGND sg13g2_nor3_1
X_4094_ net686 VGND VPWR net939 _0048_ clknet_leaf_46_clk_regs sg13g2_dfrbpq_1
XFILLER_49_891 VPWR VGND sg13g2_decap_8
X_3045_ net647 VPWR _1132_ VGND net933 _1033_ sg13g2_o21ai_1
XFILLER_36_541 VPWR VGND sg13g2_decap_4
XFILLER_36_596 VPWR VGND sg13g2_fill_1
XFILLER_36_585 VPWR VGND sg13g2_decap_4
X_3947_ VGND VPWR net57 _1799_ _0390_ _1801_ sg13g2_a21oi_1
XFILLER_23_27 VPWR VGND sg13g2_fill_2
XFILLER_20_964 VPWR VGND sg13g2_decap_4
X_3878_ _1750_ net366 _0371_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_50_clk_regs clknet_3_1__leaf_clk_regs clknet_leaf_50_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2829_ _1002_ net838 _0479_ _0522_ VPWR VGND sg13g2_and3_1
XFILLER_24_1026 VPWR VGND sg13g2_fill_2
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_47_817 VPWR VGND sg13g2_decap_8
XFILLER_48_68 VPWR VGND sg13g2_fill_1
XFILLER_27_563 VPWR VGND sg13g2_decap_4
XFILLER_14_213 VPWR VGND sg13g2_fill_1
XFILLER_27_585 VPWR VGND sg13g2_decap_4
XFILLER_15_747 VPWR VGND sg13g2_decap_4
XFILLER_42_544 VPWR VGND sg13g2_fill_1
XFILLER_7_979 VPWR VGND sg13g2_decap_8
XFILLER_9_1009 VPWR VGND sg13g2_decap_8
XFILLER_36_8 VPWR VGND sg13g2_decap_4
XFILLER_49_132 VPWR VGND sg13g2_fill_1
XFILLER_38_828 VPWR VGND sg13g2_fill_1
XFILLER_46_883 VPWR VGND sg13g2_decap_8
X_3801_ net592 _1692_ net1005 _1696_ VPWR VGND sg13g2_nand3_1
XFILLER_14_791 VPWR VGND sg13g2_fill_2
XFILLER_9_250 VPWR VGND sg13g2_fill_1
X_3732_ VPWR VGND _1499_ net627 _1633_ net637 _1634_ _1626_ sg13g2_a221oi_1
X_3663_ net777 VPWR _1567_ VGND _1565_ _1566_ sg13g2_o21ai_1
X_2614_ _0831_ net589 net471 net591 net849 VPWR VGND sg13g2_a22oi_1
X_3594_ net777 net774 _1500_ VPWR VGND sg13g2_nor2b_2
X_2545_ _0769_ u_usb_cdc.u_ctrl_endp.req_q\[6\] _0772_ VPWR VGND sg13g2_nor2b_1
X_2476_ _0701_ _0702_ _0699_ _0704_ VPWR VGND _0703_ sg13g2_nand4_1
X_4215_ net668 VGND VPWR net464 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[61\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_4146_ net661 VGND VPWR _0075_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_2
XFILLER_29_817 VPWR VGND sg13g2_fill_2
X_4077_ _1897_ net404 _1898_ VPWR VGND sg13g2_xor2_1
X_3028_ _1122_ VPWR _0150_ VGND _1087_ _1098_ sg13g2_o21ai_1
XFILLER_12_728 VPWR VGND sg13g2_decap_4
XFILLER_11_238 VPWR VGND sg13g2_fill_1
Xclkload3 clkload3/Y clknet_leaf_21_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_8_1020 VPWR VGND sg13g2_decap_8
XFILLER_30_569 VPWR VGND sg13g2_fill_2
XFILLER_30_558 VPWR VGND sg13g2_fill_2
XFILLER_10_282 VPWR VGND sg13g2_fill_1
XFILLER_3_982 VPWR VGND sg13g2_decap_8
X_2330_ _0562_ _1924_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\]
+ net809 _1922_ VPWR VGND sg13g2_a22oi_1
XFILLER_2_470 VPWR VGND sg13g2_fill_1
X_2261_ _0493_ net967 u_usb_cdc.u_sie.data_q\[5\] VPWR VGND sg13g2_xnor2_1
X_4000_ net709 VPWR _1834_ VGND net835 _0926_ sg13g2_o21ai_1
X_2192_ net310 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[4\] _2046_ VPWR VGND sg13g2_nor2_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_37_135 VPWR VGND sg13g2_fill_1
XFILLER_38_669 VPWR VGND sg13g2_fill_1
XFILLER_45_190 VPWR VGND sg13g2_fill_1
XFILLER_14_1014 VPWR VGND sg13g2_decap_8
X_3715_ VGND VPWR net798 _1616_ _1617_ net796 sg13g2_a21oi_1
X_3646_ _1551_ _1506_ _1520_ VPWR VGND sg13g2_nand2_1
X_3577_ _0326_ net579 _0494_ net583 _1964_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_407 VPWR VGND sg13g2_decap_8
XFILLER_1_919 VPWR VGND sg13g2_decap_8
X_2528_ _0755_ _0754_ _0748_ _0753_ _0719_ VPWR VGND sg13g2_a22oi_1
Xhold15 _0390_ VPWR VGND net58 sg13g2_dlygate4sd3_1
X_2459_ u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\]
+ u_usb_cdc.configured_o VPWR VGND sg13g2_and2_1
Xhold37 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[49\] VPWR VGND
+ net80 sg13g2_dlygate4sd3_1
Xhold26 _0153_ VPWR VGND net69 sg13g2_dlygate4sd3_1
Xhold59 _0224_ VPWR VGND net102 sg13g2_dlygate4sd3_1
XFILLER_21_1018 VPWR VGND sg13g2_decap_8
Xhold48 _0127_ VPWR VGND net91 sg13g2_dlygate4sd3_1
X_4129_ net695 VGND VPWR _0019_ u_usb_cdc.u_sie.phy_state_q\[11\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_43_138 VPWR VGND sg13g2_fill_2
XFILLER_4_713 VPWR VGND sg13g2_fill_1
XFILLER_10_83 VPWR VGND sg13g2_fill_1
XFILLER_0_930 VPWR VGND sg13g2_decap_8
XFILLER_48_934 VPWR VGND sg13g2_decap_8
XFILLER_34_105 VPWR VGND sg13g2_fill_2
XFILLER_47_488 VPWR VGND sg13g2_fill_2
XFILLER_47_499 VPWR VGND sg13g2_decap_8
XFILLER_35_639 VPWR VGND sg13g2_fill_1
XFILLER_31_801 VPWR VGND sg13g2_fill_1
XFILLER_42_182 VPWR VGND sg13g2_fill_1
X_3500_ _1447_ _0653_ _1446_ VPWR VGND sg13g2_nand2_1
Xhold518 _0866_ VPWR VGND net561 sg13g2_dlygate4sd3_1
Xhold507 _0084_ VPWR VGND net550 sg13g2_dlygate4sd3_1
X_4480_ net729 VGND VPWR net229 u_usb_cdc.u_sie.rx_data\[4\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_1
Xhold529 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[1\] VPWR VGND net572 sg13g2_dlygate4sd3_1
X_3431_ _1400_ _1388_ _1401_ VPWR VGND sg13g2_nor2b_2
X_3362_ _1357_ _1355_ _1356_ _1352_ net812 VPWR VGND sg13g2_a22oi_1
X_2313_ net776 net773 _0545_ VPWR VGND sg13g2_nor2_1
X_3293_ VGND VPWR net152 net629 _1295_ net617 sg13g2_a21oi_1
X_2244_ _0476_ _0466_ _0475_ VPWR VGND sg13g2_nand2_1
XFILLER_39_967 VPWR VGND sg13g2_decap_8
XFILLER_18_0 VPWR VGND sg13g2_fill_1
X_2175_ VGND VPWR _2007_ _2025_ _0066_ _2030_ sg13g2_a21oi_1
XFILLER_34_694 VPWR VGND sg13g2_decap_4
X_3629_ net602 VPWR _1535_ VGND net187 _1523_ sg13g2_o21ai_1
XFILLER_1_727 VPWR VGND sg13g2_decap_8
Xoutput16 net16 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput27 net27 usb_dn_en_o VPWR VGND sg13g2_buf_1
XFILLER_49_709 VPWR VGND sg13g2_decap_8
XFILLER_5_1012 VPWR VGND sg13g2_decap_8
XFILLER_45_904 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_5_clk_regs clknet_3_0__leaf_clk_regs clknet_leaf_5_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_40_642 VPWR VGND sg13g2_fill_1
XFILLER_39_208 VPWR VGND sg13g2_fill_1
XFILLER_48_731 VPWR VGND sg13g2_decap_8
XFILLER_44_970 VPWR VGND sg13g2_decap_8
X_3980_ _1818_ VPWR _0406_ VGND _1952_ net613 sg13g2_o21ai_1
X_2931_ _1072_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net644 VPWR VGND sg13g2_nand2_1
Xclkbuf_0_clk clk delaynet_0_clk VPWR VGND sg13g2_buf_8
X_2862_ _1033_ net547 _1032_ VPWR VGND sg13g2_nand2_2
XFILLER_30_174 VPWR VGND sg13g2_fill_2
X_2793_ _0970_ _0964_ net745 _0600_ net593 VPWR VGND sg13g2_a22oi_1
XFILLER_11_1017 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_4532_ net27 net29 VPWR VGND sg13g2_buf_1
Xhold315 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[21\] VPWR
+ VGND net358 sg13g2_dlygate4sd3_1
Xhold304 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[51\] VPWR
+ VGND net347 sg13g2_dlygate4sd3_1
Xhold326 _0037_ VPWR VGND net369 sg13g2_dlygate4sd3_1
X_4463_ net726 VGND VPWR net919 u_usb_cdc.bus_reset clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
X_3414_ VGND VPWR _1913_ net578 _0265_ _1393_ sg13g2_a21oi_1
Xhold359 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[53\] VPWR
+ VGND net402 sg13g2_dlygate4sd3_1
Xhold337 _0071_ VPWR VGND net380 sg13g2_dlygate4sd3_1
Xhold348 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[9\] VPWR VGND net391 sg13g2_dlygate4sd3_1
X_4394_ net698 VGND VPWR net401 u_usb_cdc.u_sie.in_byte_q\[3\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_1
Xfanout806 net811 net806 VPWR VGND sg13g2_buf_8
X_3345_ _1340_ VPWR _1341_ VGND net819 net255 sg13g2_o21ai_1
Xfanout839 u_usb_cdc.u_sie.phy_state_q\[9\] net839 VPWR VGND sg13g2_buf_1
Xfanout817 net1051 net817 VPWR VGND sg13g2_buf_8
Xfanout828 net268 net828 VPWR VGND sg13g2_buf_8
X_3276_ _1279_ net770 net951 VPWR VGND sg13g2_nand2_1
X_2227_ _0459_ net763 net762 VPWR VGND sg13g2_xnor2_1
XFILLER_38_241 VPWR VGND sg13g2_fill_2
X_2158_ VGND VPWR _2014_ u_usb_cdc.endp\[2\] u_usb_cdc.endp\[3\] sg13g2_or2_1
X_2089_ VPWR _1946_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] VGND sg13g2_inv_1
XFILLER_34_491 VPWR VGND sg13g2_decap_8
XFILLER_22_675 VPWR VGND sg13g2_fill_2
XFILLER_6_819 VPWR VGND sg13g2_fill_2
XFILLER_1_568 VPWR VGND sg13g2_decap_4
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_27_1024 VPWR VGND sg13g2_decap_4
XFILLER_49_506 VPWR VGND sg13g2_decap_8
XFILLER_45_712 VPWR VGND sg13g2_decap_8
XFILLER_44_200 VPWR VGND sg13g2_fill_1
XFILLER_45_745 VPWR VGND sg13g2_decap_8
XFILLER_44_233 VPWR VGND sg13g2_decap_4
XFILLER_26_981 VPWR VGND sg13g2_decap_8
XFILLER_41_984 VPWR VGND sg13g2_decap_8
XFILLER_12_185 VPWR VGND sg13g2_fill_2
XFILLER_5_841 VPWR VGND sg13g2_fill_1
XFILLER_4_362 VPWR VGND sg13g2_fill_2
X_3130_ net358 net633 _1187_ VPWR VGND sg13g2_nor2_1
X_3061_ net829 net826 _1139_ VPWR VGND sg13g2_nor2_1
XFILLER_48_550 VPWR VGND sg13g2_decap_8
XFILLER_48_572 VPWR VGND sg13g2_decap_8
X_3963_ VGND VPWR _1944_ _2040_ _0397_ net557 sg13g2_a21oi_1
X_2914_ _1060_ net644 VPWR VGND net618 sg13g2_nand2b_2
X_3894_ VGND VPWR _2004_ _1763_ _0375_ _1762_ sg13g2_a21oi_1
X_2845_ net833 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\] net977
+ _1016_ VPWR VGND sg13g2_nand3_1
Xhold101 _0200_ VPWR VGND net144 sg13g2_dlygate4sd3_1
X_2776_ _0953_ VPWR _0954_ VGND net769 _1987_ sg13g2_o21ai_1
X_4515_ net681 VGND VPWR _0427_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\]
+ clknet_leaf_20_clk_regs sg13g2_dfrbpq_1
Xhold123 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[70\] VPWR
+ VGND net166 sg13g2_dlygate4sd3_1
Xhold112 _0117_ VPWR VGND net155 sg13g2_dlygate4sd3_1
Xhold134 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[39\] VPWR VGND
+ net177 sg13g2_dlygate4sd3_1
Xhold156 _0118_ VPWR VGND net199 sg13g2_dlygate4sd3_1
X_4446_ net725 VGND VPWR net349 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[4\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
Xhold145 _0401_ VPWR VGND net188 sg13g2_dlygate4sd3_1
Xhold167 _0362_ VPWR VGND net210 sg13g2_dlygate4sd3_1
Xfanout603 net604 net603 VPWR VGND sg13g2_buf_8
X_4377_ net688 VGND VPWR _0305_ u_usb_cdc.endp\[2\] clknet_leaf_42_clk_regs sg13g2_dfrbpq_2
Xfanout614 _0942_ net614 VPWR VGND sg13g2_buf_8
Xhold178 _0097_ VPWR VGND net221 sg13g2_dlygate4sd3_1
Xhold189 u_usb_cdc.u_sie.rx_data\[2\] VPWR VGND net232 sg13g2_dlygate4sd3_1
X_3328_ _1325_ VPWR _1326_ VGND net823 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[4\]
+ sg13g2_o21ai_1
Xfanout658 net659 net658 VPWR VGND sg13g2_buf_8
Xfanout625 _2023_ net625 VPWR VGND sg13g2_buf_8
Xfanout647 _1014_ net647 VPWR VGND sg13g2_buf_8
Xfanout636 _1078_ net636 VPWR VGND sg13g2_buf_8
Xfanout669 net670 net669 VPWR VGND sg13g2_buf_8
X_3259_ net770 net830 _1265_ VPWR VGND sg13g2_nor2_1
XFILLER_39_594 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_1_332 VPWR VGND sg13g2_decap_8
XFILLER_2_855 VPWR VGND sg13g2_decap_4
Xhold690 _0060_ VPWR VGND net1009 sg13g2_dlygate4sd3_1
XFILLER_27_70 VPWR VGND sg13g2_decap_8
XFILLER_18_778 VPWR VGND sg13g2_decap_8
X_2630_ _0842_ _0455_ net593 VPWR VGND sg13g2_nand2_1
XFILLER_40_291 VPWR VGND sg13g2_decap_8
XFILLER_9_487 VPWR VGND sg13g2_fill_1
X_2561_ _0649_ _0698_ _0749_ _0787_ VPWR VGND sg13g2_nor3_1
X_2492_ _0720_ _0717_ _0719_ VPWR VGND sg13g2_nand2_2
X_4300_ net673 VGND VPWR net373 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[62\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_4231_ net679 VGND VPWR _0160_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[1\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_2
X_4162_ net680 VGND VPWR net83 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[8\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
XFILLER_49_870 VPWR VGND sg13g2_decap_8
X_3113_ net829 net739 _1175_ VPWR VGND net830 sg13g2_nand3b_1
X_4093_ net689 VGND VPWR net487 u_usb_cdc.u_sie.out_toggle_q\[0\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_1
X_3044_ net882 _1131_ _1128_ _0157_ VPWR VGND sg13g2_mux2_1
XFILLER_36_564 VPWR VGND sg13g2_decap_8
X_3946_ VGND VPWR _1796_ _1797_ _1801_ net57 sg13g2_a21oi_1
XFILLER_11_409 VPWR VGND sg13g2_decap_8
X_3877_ VGND VPWR net741 net361 _1751_ net365 sg13g2_a21oi_1
X_2828_ net379 _1001_ _0071_ VPWR VGND sg13g2_nor2b_1
X_2759_ net748 _0943_ _0045_ VPWR VGND sg13g2_nor2_1
XFILLER_2_118 VPWR VGND sg13g2_fill_1
X_4429_ net697 VGND VPWR net999 u_usb_cdc.u_sie.pid_q\[2\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1005 VPWR VGND sg13g2_decap_8
XFILLER_48_58 VPWR VGND sg13g2_fill_1
XFILLER_27_520 VPWR VGND sg13g2_fill_2
XFILLER_27_542 VPWR VGND sg13g2_decap_8
XFILLER_27_597 VPWR VGND sg13g2_fill_2
XFILLER_42_523 VPWR VGND sg13g2_decap_8
XFILLER_31_1009 VPWR VGND sg13g2_decap_8
XFILLER_6_413 VPWR VGND sg13g2_fill_2
XFILLER_13_72 VPWR VGND sg13g2_fill_1
XFILLER_7_958 VPWR VGND sg13g2_decap_8
XFILLER_2_685 VPWR VGND sg13g2_fill_1
XFILLER_2_674 VPWR VGND sg13g2_decap_8
XFILLER_2_696 VPWR VGND sg13g2_decap_8
XFILLER_49_111 VPWR VGND sg13g2_decap_8
XFILLER_38_818 VPWR VGND sg13g2_fill_2
XFILLER_49_155 VPWR VGND sg13g2_fill_1
XFILLER_46_862 VPWR VGND sg13g2_decap_8
X_3800_ _1695_ VPWR _0349_ VGND _1913_ net600 sg13g2_o21ai_1
XFILLER_33_578 VPWR VGND sg13g2_decap_4
XFILLER_20_228 VPWR VGND sg13g2_fill_1
X_3731_ _1631_ VPWR _1633_ VGND _1539_ _1632_ sg13g2_o21ai_1
X_3662_ net788 _1506_ _1566_ VPWR VGND sg13g2_nor2_1
X_2613_ _0610_ _0829_ net742 _0830_ VPWR VGND sg13g2_nand3_1
X_3593_ net849 _0551_ _0552_ _1499_ VGND VPWR _1498_ sg13g2_nor4_2
X_2544_ VGND VPWR _0692_ _0770_ _0771_ _0769_ sg13g2_a21oi_1
XFILLER_47_1027 VPWR VGND sg13g2_fill_2
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2475_ VPWR VGND net588 _0681_ _0665_ _0635_ _0703_ _0662_ sg13g2_a221oi_1
X_4214_ net668 VGND VPWR net476 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[60\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
X_4145_ net678 VGND VPWR net548 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_q
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
XFILLER_37_851 VPWR VGND sg13g2_fill_2
X_4076_ _1897_ net350 net389 VPWR VGND sg13g2_nand2_1
X_3027_ _1122_ net123 _1118_ VPWR VGND sg13g2_nand2_1
XFILLER_11_217 VPWR VGND sg13g2_fill_1
Xclkload4 VPWR clkload4/Y clknet_leaf_34_clk_regs VGND sg13g2_inv_1
X_3929_ net353 _1786_ _1789_ VPWR VGND sg13g2_and2_1
XFILLER_42_353 VPWR VGND sg13g2_decap_4
XFILLER_42_342 VPWR VGND sg13g2_fill_2
XFILLER_43_898 VPWR VGND sg13g2_decap_8
XFILLER_3_961 VPWR VGND sg13g2_decap_8
X_2260_ _0492_ net888 u_usb_cdc.u_sie.data_q\[6\] VPWR VGND sg13g2_xnor2_1
X_2191_ _1944_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\] u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[6\]
+ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[7\] _2045_ VPWR VGND sg13g2_nor4_1
XFILLER_38_615 VPWR VGND sg13g2_decap_4
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_21_537 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_29_clk_regs clknet_3_7__leaf_clk_regs clknet_leaf_29_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3714_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[20\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[28\]
+ net804 _1616_ VPWR VGND sg13g2_mux2_1
X_3645_ net779 _0542_ _0668_ _1550_ VPWR VGND sg13g2_nor3_1
X_3576_ _0325_ net579 _1495_ _1492_ _1965_ VPWR VGND sg13g2_a22oi_1
X_2527_ _0649_ net622 _0749_ _0754_ VPWR VGND sg13g2_nor3_1
X_2458_ _0061_ _0687_ _0662_ _0679_ _2005_ VPWR VGND sg13g2_a22oi_1
Xhold38 _0132_ VPWR VGND net81 sg13g2_dlygate4sd3_1
Xhold16 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[43\] VPWR VGND
+ net59 sg13g2_dlygate4sd3_1
Xhold27 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[46\] VPWR VGND
+ net70 sg13g2_dlygate4sd3_1
X_2389_ VGND VPWR _0620_ net590 _0615_ sg13g2_or2_1
Xhold49 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[64\] VPWR VGND
+ net92 sg13g2_dlygate4sd3_1
X_4128_ net703 VGND VPWR _0018_ u_usb_cdc.u_sie.phy_state_q\[10\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
X_4059_ _0922_ net937 _1885_ VPWR VGND sg13g2_xor2_1
XFILLER_25_821 VPWR VGND sg13g2_fill_1
XFILLER_12_504 VPWR VGND sg13g2_decap_8
XFILLER_12_515 VPWR VGND sg13g2_fill_1
Xclkbuf_regs_0_clk clk clk_regs VPWR VGND sg13g2_buf_8
XFILLER_48_913 VPWR VGND sg13g2_decap_8
XFILLER_0_986 VPWR VGND sg13g2_decap_8
XFILLER_19_158 VPWR VGND sg13g2_fill_1
XFILLER_16_843 VPWR VGND sg13g2_fill_2
XFILLER_16_887 VPWR VGND sg13g2_decap_8
XFILLER_35_81 VPWR VGND sg13g2_fill_2
Xhold508 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq
+ VPWR VGND net551 sg13g2_dlygate4sd3_1
X_3430_ _1398_ _1399_ _1400_ VPWR VGND sg13g2_nor2_1
Xhold519 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] VPWR VGND net562 sg13g2_dlygate4sd3_1
X_3361_ VGND VPWR net824 _2002_ _1356_ _1286_ sg13g2_a21oi_1
XFILLER_44_1019 VPWR VGND sg13g2_decap_8
X_2312_ net780 _0543_ _0544_ VPWR VGND sg13g2_nor2_1
X_3292_ net819 _1983_ _1288_ _1294_ VPWR VGND sg13g2_nor3_2
X_2243_ _0475_ u_usb_cdc.u_sie.data_q\[4\] _0468_ VPWR VGND sg13g2_xnor2_1
X_2174_ net643 net873 _2030_ VPWR VGND sg13g2_nor2_1
XFILLER_25_139 VPWR VGND sg13g2_fill_1
XFILLER_33_194 VPWR VGND sg13g2_fill_1
X_3628_ VPWR VGND net637 net627 _1533_ _1499_ _1534_ _1522_ sg13g2_a221oi_1
Xoutput28 net28 usb_dn_tx_o VPWR VGND sg13g2_buf_1
XFILLER_1_706 VPWR VGND sg13g2_decap_8
Xoutput17 net17 uio_out[6] VPWR VGND sg13g2_buf_1
X_3559_ _1484_ net376 net327 VPWR VGND sg13g2_xnor2_1
XFILLER_0_238 VPWR VGND sg13g2_decap_4
XFILLER_17_618 VPWR VGND sg13g2_fill_2
XFILLER_12_367 VPWR VGND sg13g2_fill_2
XFILLER_8_349 VPWR VGND sg13g2_fill_1
XFILLER_0_783 VPWR VGND sg13g2_decap_8
XFILLER_48_710 VPWR VGND sg13g2_decap_8
XFILLER_48_787 VPWR VGND sg13g2_decap_8
X_2930_ _1071_ net72 _1060_ VPWR VGND sg13g2_nand2_1
XFILLER_31_654 VPWR VGND sg13g2_fill_1
XFILLER_31_676 VPWR VGND sg13g2_decap_8
X_2861_ VGND VPWR _1032_ _1031_ net716 sg13g2_or2_1
X_2792_ VGND VPWR net840 _0513_ _0969_ _0968_ sg13g2_a21oi_1
X_4531_ u_usb_cdc.configured_o net17 VPWR VGND sg13g2_buf_8
X_4462_ net735 VGND VPWR net58 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[2\] clknet_leaf_27_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_7_393 VPWR VGND sg13g2_fill_2
Xhold316 _1187_ VPWR VGND net359 sg13g2_dlygate4sd3_1
Xhold305 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[4\] VPWR VGND net348 sg13g2_dlygate4sd3_1
X_3413_ net545 net578 _1393_ VPWR VGND sg13g2_nor2_1
Xhold338 u_usb_cdc.u_sie.addr_q\[5\] VPWR VGND net381 sg13g2_dlygate4sd3_1
Xhold327 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[31\] VPWR
+ VGND net370 sg13g2_dlygate4sd3_1
Xhold349 _0379_ VPWR VGND net392 sg13g2_dlygate4sd3_1
X_4393_ net697 VGND VPWR net322 u_usb_cdc.u_sie.in_byte_q\[2\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_1
Xfanout807 net811 net807 VPWR VGND sg13g2_buf_8
X_3344_ VGND VPWR net819 _2000_ _1340_ net815 sg13g2_a21oi_1
Xfanout818 net819 net818 VPWR VGND sg13g2_buf_8
Xfanout829 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\] net829
+ VPWR VGND sg13g2_buf_8
X_3275_ _1278_ _0714_ _1252_ VPWR VGND sg13g2_nand2_1
X_2226_ _0458_ _0456_ _0457_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_231 VPWR VGND sg13g2_fill_1
X_2157_ VPWR _2013_ net264 VGND sg13g2_inv_1
XFILLER_26_39 VPWR VGND sg13g2_decap_8
X_2088_ VPWR _1945_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\] VGND sg13g2_inv_1
Xclkbuf_leaf_44_clk_regs clknet_3_4__leaf_clk_regs clknet_leaf_44_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_42_16 VPWR VGND sg13g2_decap_4
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_27_1003 VPWR VGND sg13g2_decap_8
XFILLER_26_960 VPWR VGND sg13g2_decap_8
XFILLER_41_963 VPWR VGND sg13g2_decap_8
XFILLER_12_142 VPWR VGND sg13g2_fill_2
XFILLER_9_658 VPWR VGND sg13g2_fill_2
XFILLER_40_495 VPWR VGND sg13g2_decap_4
XFILLER_5_875 VPWR VGND sg13g2_decap_8
X_3060_ _1138_ VPWR _0166_ VGND _1924_ _1135_ sg13g2_o21ai_1
XFILLER_48_540 VPWR VGND sg13g2_decap_4
XFILLER_48_584 VPWR VGND sg13g2_decap_8
X_3962_ net556 _2040_ _1810_ VPWR VGND sg13g2_nor2_1
X_2913_ net834 net833 _1059_ VPWR VGND sg13g2_nor2b_2
X_3893_ net348 _1754_ net741 _1763_ VPWR VGND sg13g2_nand3_1
XFILLER_31_484 VPWR VGND sg13g2_decap_8
XFILLER_32_996 VPWR VGND sg13g2_decap_8
X_2844_ _1015_ net834 net833 VPWR VGND sg13g2_nand2_2
XFILLER_8_691 VPWR VGND sg13g2_fill_2
X_2775_ _0953_ net769 u_usb_cdc.u_sie.out_toggle_q\[1\] VPWR VGND sg13g2_nand2_1
X_4514_ net705 VGND VPWR net165 u_usb_cdc.u_sie.in_zlp_q\[0\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_1
Xhold102 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[25\] VPWR
+ VGND net145 sg13g2_dlygate4sd3_1
Xhold124 _0237_ VPWR VGND net167 sg13g2_dlygate4sd3_1
Xhold113 u_usb_cdc.u_sie.delay_cnt_q\[2\] VPWR VGND net156 sg13g2_dlygate4sd3_1
Xhold135 _0122_ VPWR VGND net178 sg13g2_dlygate4sd3_1
Xhold168 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[59\] VPWR
+ VGND net211 sg13g2_dlygate4sd3_1
Xhold146 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[37\] VPWR
+ VGND net189 sg13g2_dlygate4sd3_1
Xhold157 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[65\] VPWR VGND
+ net200 sg13g2_dlygate4sd3_1
X_4445_ net725 VGND VPWR net983 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[3\] clknet_leaf_19_clk_regs
+ sg13g2_dfrbpq_1
X_4376_ net687 VGND VPWR _0304_ u_usb_cdc.endp\[1\] clknet_leaf_42_clk_regs sg13g2_dfrbpq_2
Xfanout604 _1232_ net604 VPWR VGND sg13g2_buf_8
Xhold179 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[14\] VPWR
+ VGND net222 sg13g2_dlygate4sd3_1
Xfanout615 _1746_ net615 VPWR VGND sg13g2_buf_8
X_3327_ _1325_ net823 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[12\]
+ VPWR VGND sg13g2_nand2b_1
Xfanout648 net651 net648 VPWR VGND sg13g2_buf_8
Xfanout626 _2020_ net626 VPWR VGND sg13g2_buf_8
Xfanout637 net638 net637 VPWR VGND sg13g2_buf_2
Xfanout659 net671 net659 VPWR VGND sg13g2_buf_8
X_3258_ _1264_ _1263_ VPWR VGND _1249_ sg13g2_nand2b_2
XFILLER_39_562 VPWR VGND sg13g2_decap_4
X_3189_ _1220_ VPWR _0213_ VGND net711 _1172_ sg13g2_o21ai_1
X_2209_ _0441_ net838 net750 VPWR VGND sg13g2_nand2b_1
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_41_204 VPWR VGND sg13g2_fill_2
XFILLER_23_985 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_fill_2
XFILLER_22_484 VPWR VGND sg13g2_fill_2
Xhold680 _0357_ VPWR VGND net999 sg13g2_dlygate4sd3_1
Xhold691 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ VPWR VGND net1010 sg13g2_dlygate4sd3_1
XFILLER_1_388 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_4
XFILLER_17_245 VPWR VGND sg13g2_fill_1
XFILLER_17_223 VPWR VGND sg13g2_fill_1
XFILLER_45_598 VPWR VGND sg13g2_fill_2
XFILLER_9_400 VPWR VGND sg13g2_fill_2
X_2560_ _0786_ _0641_ _0694_ VPWR VGND sg13g2_nand2_1
X_2491_ net787 net715 _0635_ _0719_ VGND VPWR _0675_ sg13g2_nor4_2
X_4230_ net678 VGND VPWR net978 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[0\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_2
X_4161_ net678 VGND VPWR net870 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[7\]
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
X_3112_ _1173_ VPWR _0182_ VGND u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[2\]
+ _1174_ sg13g2_o21ai_1
X_4092_ _0053_ net27 VPWR VGND sg13g2_buf_1
X_3043_ _1021_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] _1031_
+ _1131_ VPWR VGND sg13g2_mux2_1
XFILLER_36_554 VPWR VGND sg13g2_fill_1
X_3945_ _1799_ net424 _0389_ VPWR VGND sg13g2_nor2_1
XFILLER_17_1013 VPWR VGND sg13g2_decap_8
XFILLER_23_18 VPWR VGND sg13g2_fill_1
XFILLER_31_270 VPWR VGND sg13g2_fill_2
X_3876_ net716 _1749_ _1750_ VPWR VGND sg13g2_nor2_1
X_2827_ _0995_ VPWR _1001_ VGND net851 _1000_ sg13g2_o21ai_1
X_2758_ net450 net614 _0943_ VPWR VGND sg13g2_nor2b_1
X_2689_ _0888_ _0889_ _0885_ _0890_ VPWR VGND sg13g2_nand3_1
X_4428_ net697 VGND VPWR net945 u_usb_cdc.u_sie.pid_q\[1\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_2
X_4359_ net686 VGND VPWR _0287_ u_usb_cdc.u_ctrl_endp.in_dir_q clknet_leaf_47_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_922 VPWR VGND sg13g2_decap_4
XFILLER_23_782 VPWR VGND sg13g2_decap_8
XFILLER_6_469 VPWR VGND sg13g2_fill_2
XFILLER_6_458 VPWR VGND sg13g2_decap_8
XFILLER_38_808 VPWR VGND sg13g2_decap_4
XFILLER_46_841 VPWR VGND sg13g2_decap_8
XFILLER_45_362 VPWR VGND sg13g2_fill_2
X_3730_ _1632_ _1520_ _1607_ VPWR VGND sg13g2_nand2_1
X_3661_ VGND VPWR _0533_ _0541_ _1565_ net780 sg13g2_a21oi_1
X_2612_ _1927_ _0595_ _0615_ _0829_ VPWR VGND sg13g2_nor3_1
X_3592_ _1498_ _0549_ net637 VPWR VGND sg13g2_nand2b_1
X_2543_ VGND VPWR net764 _1936_ _0770_ u_usb_cdc.u_ctrl_endp.rec_q\[1\] sg13g2_a21oi_1
XFILLER_47_1006 VPWR VGND sg13g2_decap_8
XFILLER_5_480 VPWR VGND sg13g2_decap_8
X_2474_ _0702_ _0663_ net623 VPWR VGND sg13g2_nand2_1
X_4213_ net667 VGND VPWR net468 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[59\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
X_4144_ net702 VGND VPWR net300 _0054_ clknet_leaf_37_clk_regs sg13g2_dfrbpq_1
XFILLER_18_29 VPWR VGND sg13g2_fill_2
X_4075_ _1896_ net404 net718 VPWR VGND sg13g2_nand2_1
X_3026_ _1121_ VPWR _0149_ VGND _1085_ _1098_ sg13g2_o21ai_1
Xclkload5 clknet_leaf_27_clk_regs clkload5/Y VPWR VGND sg13g2_inv_4
X_3928_ _1788_ net714 net353 VPWR VGND sg13g2_nand2_1
XFILLER_20_785 VPWR VGND sg13g2_decap_4
XFILLER_30_1010 VPWR VGND sg13g2_decap_8
X_3859_ _1736_ VPWR _0367_ VGND _1952_ net595 sg13g2_o21ai_1
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_47_649 VPWR VGND sg13g2_decap_8
XFILLER_15_502 VPWR VGND sg13g2_fill_1
XFILLER_43_855 VPWR VGND sg13g2_fill_2
XFILLER_42_376 VPWR VGND sg13g2_fill_2
XFILLER_24_61 VPWR VGND sg13g2_fill_1
XFILLER_23_590 VPWR VGND sg13g2_fill_1
XFILLER_11_763 VPWR VGND sg13g2_fill_2
X_2190_ _2044_ net961 _2042_ VPWR VGND sg13g2_nand2_1
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_4
XFILLER_14_590 VPWR VGND sg13g2_fill_1
XFILLER_21_549 VPWR VGND sg13g2_fill_2
X_3713_ VGND VPWR net804 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[12\]
+ _1615_ _1614_ sg13g2_a21oi_1
X_3644_ _1547_ _1548_ _1542_ _1549_ VPWR VGND sg13g2_nand3_1
XFILLER_20_19 VPWR VGND sg13g2_fill_1
X_3575_ _1495_ _0492_ _0501_ VPWR VGND sg13g2_xnor2_1
X_2526_ _0751_ _0752_ _0750_ _0753_ VPWR VGND sg13g2_nand3_1
X_2457_ net759 net758 _0683_ _0686_ _0687_ VPWR VGND sg13g2_nor4_1
Xhold17 _0126_ VPWR VGND net60 sg13g2_dlygate4sd3_1
Xhold28 _0129_ VPWR VGND net71 sg13g2_dlygate4sd3_1
Xhold39 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[8\] VPWR VGND
+ net82 sg13g2_dlygate4sd3_1
X_2388_ _0619_ net590 VPWR VGND sg13g2_inv_2
X_4127_ net687 VGND VPWR net505 u_usb_cdc.u_sie.phy_state_q\[9\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_126 VPWR VGND sg13g2_fill_1
XFILLER_29_649 VPWR VGND sg13g2_fill_1
X_4058_ net643 _1010_ _1884_ VPWR VGND sg13g2_nor2_1
XFILLER_44_619 VPWR VGND sg13g2_fill_1
X_3009_ _1116_ net150 _1108_ VPWR VGND sg13g2_nand2_1
XFILLER_40_869 VPWR VGND sg13g2_fill_1
XFILLER_40_858 VPWR VGND sg13g2_fill_2
XFILLER_0_965 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_fill_2
XFILLER_48_969 VPWR VGND sg13g2_decap_8
XFILLER_19_83 VPWR VGND sg13g2_fill_2
XFILLER_19_61 VPWR VGND sg13g2_decap_8
XFILLER_47_468 VPWR VGND sg13g2_fill_2
XFILLER_47_457 VPWR VGND sg13g2_decap_8
XFILLER_34_107 VPWR VGND sg13g2_fill_1
XFILLER_28_682 VPWR VGND sg13g2_fill_1
XFILLER_37_1027 VPWR VGND sg13g2_fill_2
Xhold509 _1907_ VPWR VGND net552 sg13g2_dlygate4sd3_1
X_3360_ VGND VPWR _1355_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[23\]
+ net824 sg13g2_or2_1
X_2311_ net788 net791 _0543_ VPWR VGND net784 sg13g2_nand3b_1
X_3291_ VPWR VGND _1289_ _1292_ _1287_ net812 _1293_ _1285_ sg13g2_a221oi_1
XFILLER_32_4 VPWR VGND sg13g2_fill_2
X_2242_ _0471_ _0472_ u_usb_cdc.u_sie.data_q\[7\] _0474_ VPWR VGND sg13g2_mux2_1
X_2173_ _2029_ _2028_ net872 net709 net835 VPWR VGND sg13g2_a22oi_1
XFILLER_34_674 VPWR VGND sg13g2_decap_8
XFILLER_22_858 VPWR VGND sg13g2_fill_1
X_3627_ _1525_ VPWR _1533_ VGND net795 _1532_ sg13g2_o21ai_1
Xoutput29 net29 usb_dp_en_o VPWR VGND sg13g2_buf_1
Xoutput18 net18 uio_out[7] VPWR VGND sg13g2_buf_1
X_3558_ _1483_ net376 net598 VPWR VGND sg13g2_nand2_1
X_2509_ net721 _0719_ net764 _0736_ VPWR VGND sg13g2_nand3_1
X_3489_ _1436_ _1438_ net588 _1439_ VPWR VGND sg13g2_nand3_1
XFILLER_45_939 VPWR VGND sg13g2_decap_8
XFILLER_16_129 VPWR VGND sg13g2_fill_2
XFILLER_25_652 VPWR VGND sg13g2_fill_2
XFILLER_40_677 VPWR VGND sg13g2_fill_1
XFILLER_0_762 VPWR VGND sg13g2_decap_8
XFILLER_48_766 VPWR VGND sg13g2_decap_8
XFILLER_29_980 VPWR VGND sg13g2_decap_8
X_2860_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_valid_qq
+ VPWR _1031_ VGND _1022_ _1030_ sg13g2_o21ai_1
X_2791_ _0968_ _0438_ _0967_ VPWR VGND sg13g2_nand2_1
XFILLER_8_862 VPWR VGND sg13g2_decap_8
XFILLER_30_198 VPWR VGND sg13g2_fill_2
X_4530_ u_usb_cdc.in_ready_o[0] net16 VPWR VGND sg13g2_buf_1
X_4461_ net735 VGND VPWR net425 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\] clknet_leaf_26_clk_regs
+ sg13g2_dfrbpq_1
Xhold317 _0188_ VPWR VGND net360 sg13g2_dlygate4sd3_1
Xhold306 _0374_ VPWR VGND net349 sg13g2_dlygate4sd3_1
X_3412_ VGND VPWR net721 _1390_ _0264_ _1392_ sg13g2_a21oi_1
Xhold339 _0311_ VPWR VGND net382 sg13g2_dlygate4sd3_1
Xhold328 _0198_ VPWR VGND net371 sg13g2_dlygate4sd3_1
X_4392_ net703 VGND VPWR net377 u_usb_cdc.u_sie.in_byte_q\[1\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_2
X_3343_ VGND VPWR _2011_ net616 _0248_ _1339_ sg13g2_a21oi_1
Xfanout819 net820 net819 VPWR VGND sg13g2_buf_2
Xfanout808 net811 net808 VPWR VGND sg13g2_buf_2
X_3274_ _1264_ net828 _1277_ _0241_ VPWR VGND sg13g2_a21o_1
X_2225_ net767 net760 _0457_ VPWR VGND sg13g2_xor2_1
XFILLER_27_906 VPWR VGND sg13g2_fill_1
XFILLER_38_243 VPWR VGND sg13g2_fill_1
X_2156_ VPWR _2012_ net294 VGND sg13g2_inv_1
XFILLER_26_18 VPWR VGND sg13g2_decap_8
X_2087_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\] _1944_ VPWR VGND sg13g2_inv_4
XFILLER_35_983 VPWR VGND sg13g2_decap_8
XFILLER_22_611 VPWR VGND sg13g2_decap_8
XFILLER_22_644 VPWR VGND sg13g2_decap_8
XFILLER_22_677 VPWR VGND sg13g2_fill_1
XFILLER_22_655 VPWR VGND sg13g2_fill_1
XFILLER_10_828 VPWR VGND sg13g2_fill_1
XFILLER_22_688 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk_regs clknet_3_2__leaf_clk_regs clknet_leaf_13_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2989_ _1105_ VPWR _0128_ VGND _1054_ net611 sg13g2_o21ai_1
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_18_917 VPWR VGND sg13g2_fill_1
XFILLER_29_276 VPWR VGND sg13g2_decap_8
XFILLER_26_950 VPWR VGND sg13g2_fill_1
XFILLER_44_279 VPWR VGND sg13g2_decap_4
XFILLER_41_942 VPWR VGND sg13g2_decap_8
XFILLER_34_1008 VPWR VGND sg13g2_decap_8
XFILLER_5_865 VPWR VGND sg13g2_decap_4
XFILLER_4_364 VPWR VGND sg13g2_fill_1
XFILLER_48_530 VPWR VGND sg13g2_fill_1
X_3961_ VGND VPWR _1943_ _2040_ _0396_ net554 sg13g2_a21oi_1
XFILLER_35_257 VPWR VGND sg13g2_fill_1
X_2912_ _1057_ VPWR _0098_ VGND net620 _1058_ sg13g2_o21ai_1
XFILLER_32_975 VPWR VGND sg13g2_decap_8
X_3892_ net713 _1761_ _1762_ VPWR VGND sg13g2_nor2_1
X_2843_ _1014_ net933 net10 VPWR VGND sg13g2_nand2_1
X_2774_ _0522_ _0949_ _0512_ _0952_ VPWR VGND _0951_ sg13g2_nand4_1
X_4513_ net705 VGND VPWR net85 u_usb_cdc.u_sie.in_zlp_q\[1\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_1
Xhold103 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[41\] VPWR
+ VGND net146 sg13g2_dlygate4sd3_1
Xhold125 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[17\] VPWR VGND
+ net168 sg13g2_dlygate4sd3_1
Xhold114 _0318_ VPWR VGND net157 sg13g2_dlygate4sd3_1
Xhold147 _0204_ VPWR VGND net190 sg13g2_dlygate4sd3_1
Xhold136 u_usb_cdc.u_ctrl_endp.dev_state_q\[1\] VPWR VGND net179 sg13g2_dlygate4sd3_1
Xhold158 _0148_ VPWR VGND net201 sg13g2_dlygate4sd3_1
X_4444_ net725 VGND VPWR net337 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[2\] clknet_leaf_19_clk_regs
+ sg13g2_dfrbpq_1
X_4375_ net677 VGND VPWR _0303_ u_usb_cdc.endp\[0\] clknet_leaf_48_clk_regs sg13g2_dfrbpq_2
Xhold169 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[39\] VPWR
+ VGND net212 sg13g2_dlygate4sd3_1
Xfanout605 net607 net605 VPWR VGND sg13g2_buf_8
X_3326_ net823 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[36\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[44\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[52\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[60\] net816 _1324_
+ VPWR VGND sg13g2_mux4_1
Xfanout649 net651 net649 VPWR VGND sg13g2_buf_8
Xfanout616 net617 net616 VPWR VGND sg13g2_buf_8
Xfanout627 _1524_ net627 VPWR VGND sg13g2_buf_8
Xfanout638 net639 net638 VPWR VGND sg13g2_buf_8
X_3257_ _0714_ VPWR _1263_ VGND net770 _1262_ sg13g2_o21ai_1
XFILLER_39_530 VPWR VGND sg13g2_decap_4
X_3188_ _1220_ net234 _1213_ VPWR VGND sg13g2_nand2_1
XFILLER_2_1017 VPWR VGND sg13g2_decap_8
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
X_2208_ _0440_ net745 _0438_ VPWR VGND sg13g2_nand2_1
X_2139_ VPWR _1995_ net290 VGND sg13g2_inv_1
XFILLER_35_780 VPWR VGND sg13g2_fill_2
XFILLER_23_975 VPWR VGND sg13g2_fill_1
Xhold670 u_usb_cdc.u_sie.data_q\[5\] VPWR VGND net989 sg13g2_dlygate4sd3_1
Xhold681 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ VPWR VGND net1000 sg13g2_dlygate4sd3_1
XFILLER_1_367 VPWR VGND sg13g2_decap_8
Xhold692 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[0\] VPWR VGND net1011 sg13g2_dlygate4sd3_1
XFILLER_49_316 VPWR VGND sg13g2_fill_1
XFILLER_9_456 VPWR VGND sg13g2_fill_2
XFILLER_5_651 VPWR VGND sg13g2_decap_8
X_2490_ net789 _0539_ _0718_ VPWR VGND sg13g2_nor2_1
X_4160_ net664 VGND VPWR net527 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[6\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_3111_ net832 _1159_ net757 _1174_ VPWR VGND sg13g2_nand3_1
X_4091_ VPWR _0428_ net552 VGND sg13g2_inv_1
X_3042_ net862 _1130_ _1128_ _0156_ VPWR VGND sg13g2_mux2_1
XFILLER_36_511 VPWR VGND sg13g2_fill_1
X_3944_ VGND VPWR u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] _1796_ _1800_ net423
+ sg13g2_a21oi_1
X_3875_ VGND VPWR net361 net365 _1749_ _1745_ sg13g2_a21oi_1
X_2826_ u_usb_cdc.u_ctrl_endp.endp_q\[0\] u_usb_cdc.u_ctrl_endp.endp_q\[2\] u_usb_cdc.u_ctrl_endp.endp_q\[3\]
+ _0999_ _1000_ VPWR VGND sg13g2_nor4_1
X_2757_ VGND VPWR _0942_ _0908_ net707 sg13g2_or2_1
X_2688_ _2036_ _0884_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] _0889_ VPWR VGND
+ sg13g2_nand3_1
X_4427_ net697 VGND VPWR net912 u_usb_cdc.u_sie.pid_q\[0\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
X_4358_ net686 VGND VPWR net493 u_usb_cdc.u_ctrl_endp.class_q clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_48_49 VPWR VGND sg13g2_decap_8
X_4289_ net672 VGND VPWR _0218_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[51\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_3309_ VGND VPWR net821 _1995_ _1309_ _1286_ sg13g2_a21oi_1
XFILLER_27_522 VPWR VGND sg13g2_fill_1
XFILLER_27_599 VPWR VGND sg13g2_fill_1
XFILLER_11_901 VPWR VGND sg13g2_fill_1
XFILLER_10_433 VPWR VGND sg13g2_decap_4
XFILLER_46_820 VPWR VGND sg13g2_fill_2
XFILLER_46_897 VPWR VGND sg13g2_decap_8
XFILLER_14_772 VPWR VGND sg13g2_fill_1
XFILLER_13_271 VPWR VGND sg13g2_fill_1
XFILLER_9_275 VPWR VGND sg13g2_decap_4
X_3660_ _0762_ net781 _0544_ _1564_ VPWR VGND sg13g2_a21o_1
X_2611_ _0827_ _0828_ _0632_ _0012_ VPWR VGND sg13g2_nand3_1
X_3591_ _1497_ net488 net597 VPWR VGND sg13g2_nand2_1
X_2542_ _0683_ _0767_ _0768_ _0769_ VPWR VGND sg13g2_nor3_1
XFILLER_6_993 VPWR VGND sg13g2_decap_8
X_2473_ net623 VPWR _0701_ VGND _0637_ _0641_ sg13g2_o21ai_1
X_4212_ net666 VGND VPWR net470 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[58\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_4143_ net703 VGND VPWR _0038_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_2
X_4074_ _1894_ VPWR _0423_ VGND _1892_ _1895_ sg13g2_o21ai_1
XFILLER_37_820 VPWR VGND sg13g2_fill_1
X_3025_ _1121_ net109 _1118_ VPWR VGND sg13g2_nand2_1
XFILLER_20_731 VPWR VGND sg13g2_decap_8
XFILLER_20_742 VPWR VGND sg13g2_fill_1
X_3927_ _1785_ VPWR _0384_ VGND _1786_ _1787_ sg13g2_o21ai_1
X_3858_ _0899_ _1729_ net496 _1736_ VPWR VGND sg13g2_nand3_1
X_2809_ net768 u_usb_cdc.endp\[1\] net406 _2014_ _0985_ VPWR VGND sg13g2_nor4_1
X_3789_ VPWR _1688_ _1687_ VGND sg13g2_inv_1
XFILLER_47_606 VPWR VGND sg13g2_decap_8
XFILLER_47_628 VPWR VGND sg13g2_decap_8
XFILLER_28_897 VPWR VGND sg13g2_fill_2
XFILLER_23_580 VPWR VGND sg13g2_fill_1
XFILLER_10_241 VPWR VGND sg13g2_fill_2
XFILLER_6_256 VPWR VGND sg13g2_fill_1
XFILLER_3_996 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_45_171 VPWR VGND sg13g2_fill_1
XFILLER_46_683 VPWR VGND sg13g2_decap_8
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_3712_ net804 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[4\] _1614_
+ VPWR VGND sg13g2_nor2b_1
X_3643_ VGND VPWR _1500_ _1545_ _1548_ _1513_ sg13g2_a21oi_1
X_3574_ _0324_ net580 _0497_ net584 _1963_ VPWR VGND sg13g2_a22oi_1
X_2525_ u_usb_cdc.u_ctrl_endp.req_q\[3\] u_usb_cdc.u_ctrl_endp.req_q\[10\] u_usb_cdc.u_ctrl_endp.req_q\[9\]
+ _0752_ VPWR VGND sg13g2_nor3_1
X_2456_ _0686_ _0634_ _0685_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_38_clk_regs clknet_3_5__leaf_clk_regs clknet_leaf_38_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_29_18 VPWR VGND sg13g2_decap_8
Xhold29 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[21\] VPWR VGND
+ net72 sg13g2_dlygate4sd3_1
Xhold18 u_usb_cdc.clk_cnt_q\[1\] VPWR VGND net61 sg13g2_dlygate4sd3_1
X_4126_ net695 VGND VPWR _0027_ u_usb_cdc.u_sie.phy_state_q\[8\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
X_2387_ net743 VPWR _0618_ VGND _0594_ _0606_ sg13g2_o21ai_1
XFILLER_29_628 VPWR VGND sg13g2_decap_8
XFILLER_28_116 VPWR VGND sg13g2_fill_1
X_4057_ VGND VPWR net308 _2023_ _0418_ _1883_ sg13g2_a21oi_1
X_3008_ _1115_ VPWR _0137_ VGND _1074_ net611 sg13g2_o21ai_1
XFILLER_36_193 VPWR VGND sg13g2_fill_2
XFILLER_3_204 VPWR VGND sg13g2_fill_2
XFILLER_0_944 VPWR VGND sg13g2_decap_8
XFILLER_48_948 VPWR VGND sg13g2_decap_8
XFILLER_19_138 VPWR VGND sg13g2_fill_2
XFILLER_47_425 VPWR VGND sg13g2_decap_8
XFILLER_37_1006 VPWR VGND sg13g2_decap_8
XFILLER_31_815 VPWR VGND sg13g2_fill_2
XFILLER_7_543 VPWR VGND sg13g2_decap_4
XFILLER_7_587 VPWR VGND sg13g2_decap_4
XFILLER_3_771 VPWR VGND sg13g2_fill_2
X_3290_ _1286_ _1290_ _1291_ _1292_ VPWR VGND sg13g2_nor3_1
X_2310_ net784 _0541_ _0542_ VPWR VGND sg13g2_nor2_1
X_2241_ _0473_ _0471_ _0472_ _0466_ _1960_ VPWR VGND sg13g2_a22oi_1
XFILLER_25_4 VPWR VGND sg13g2_decap_8
X_2172_ net626 _2027_ _2028_ VPWR VGND sg13g2_nor2_2
XFILLER_47_992 VPWR VGND sg13g2_decap_8
XFILLER_34_653 VPWR VGND sg13g2_decap_4
X_3626_ _1531_ VPWR _1532_ VGND net797 _1526_ sg13g2_o21ai_1
Xoutput19 net19 uo_out[0] VPWR VGND sg13g2_buf_1
X_3557_ _1482_ VPWR _0319_ VGND net327 _0867_ sg13g2_o21ai_1
X_2508_ _0735_ _0733_ _0723_ _0732_ _0690_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_218 VPWR VGND sg13g2_decap_8
X_3488_ _1929_ VPWR _1438_ VGND _0551_ _0602_ sg13g2_o21ai_1
X_2439_ VGND VPWR _0669_ net788 net791 sg13g2_or2_1
XFILLER_5_1026 VPWR VGND sg13g2_fill_2
XFILLER_45_918 VPWR VGND sg13g2_decap_8
X_4109_ net687 VGND VPWR net380 u_usb_cdc.u_sie.in_toggle_q\[2\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_38_981 VPWR VGND sg13g2_decap_8
XFILLER_0_741 VPWR VGND sg13g2_decap_8
XFILLER_43_1010 VPWR VGND sg13g2_decap_8
XFILLER_48_745 VPWR VGND sg13g2_decap_8
XFILLER_47_288 VPWR VGND sg13g2_fill_1
XFILLER_44_984 VPWR VGND sg13g2_decap_8
XFILLER_30_111 VPWR VGND sg13g2_fill_1
XFILLER_31_645 VPWR VGND sg13g2_decap_8
XFILLER_43_494 VPWR VGND sg13g2_fill_2
X_2790_ net752 _0964_ _0967_ VPWR VGND sg13g2_nor2_1
X_4460_ net735 VGND VPWR _0388_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] clknet_leaf_27_clk_regs
+ sg13g2_dfrbpq_2
Xhold307 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] VPWR VGND net350 sg13g2_dlygate4sd3_1
X_3411_ net871 net578 _1392_ VPWR VGND sg13g2_nor2_1
Xhold329 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[62\] VPWR
+ VGND net372 sg13g2_dlygate4sd3_1
X_4391_ net697 VGND VPWR net328 u_usb_cdc.u_sie.in_byte_q\[0\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_2
Xhold318 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[0\] VPWR VGND net361 sg13g2_dlygate4sd3_1
X_3342_ VPWR VGND _1983_ net617 _1338_ net226 _1339_ _1294_ sg13g2_a221oi_1
Xfanout809 net810 net809 VPWR VGND sg13g2_buf_8
X_3273_ VGND VPWR _1275_ _1276_ _1277_ _1264_ sg13g2_a21oi_1
X_2224_ u_usb_cdc.sie_out_data\[5\] net761 _0456_ VPWR VGND sg13g2_xor2_1
XFILLER_39_723 VPWR VGND sg13g2_fill_2
X_2155_ VPWR _2011_ net244 VGND sg13g2_inv_1
XFILLER_16_0 VPWR VGND sg13g2_fill_2
XFILLER_38_222 VPWR VGND sg13g2_fill_2
XFILLER_27_929 VPWR VGND sg13g2_fill_2
X_2086_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] _1943_ VPWR VGND sg13g2_inv_4
X_2988_ _1105_ net117 _1096_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_53_clk_regs clknet_3_0__leaf_clk_regs clknet_leaf_53_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3609_ _0535_ _0674_ _1515_ VPWR VGND sg13g2_nor2_1
XFILLER_45_726 VPWR VGND sg13g2_decap_4
XFILLER_26_940 VPWR VGND sg13g2_fill_1
XFILLER_45_759 VPWR VGND sg13g2_decap_8
XFILLER_41_910 VPWR VGND sg13g2_fill_2
XFILLER_16_30 VPWR VGND sg13g2_fill_2
XFILLER_26_995 VPWR VGND sg13g2_decap_8
XFILLER_9_605 VPWR VGND sg13g2_decap_4
XFILLER_40_431 VPWR VGND sg13g2_fill_1
XFILLER_41_998 VPWR VGND sg13g2_decap_8
XFILLER_4_310 VPWR VGND sg13g2_fill_2
XFILLER_0_582 VPWR VGND sg13g2_decap_8
XFILLER_35_236 VPWR VGND sg13g2_fill_2
X_3960_ net553 _2040_ _1809_ VPWR VGND sg13g2_nor2_1
X_2911_ _1058_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ _1039_ VPWR VGND sg13g2_nand2_1
XFILLER_44_781 VPWR VGND sg13g2_decap_8
X_3891_ _1745_ _1760_ _1761_ VPWR VGND sg13g2_nor2_1
X_2842_ _1007_ VPWR _0073_ VGND _1012_ _1013_ sg13g2_o21ai_1
X_2773_ VGND VPWR _0951_ net839 net840 sg13g2_or2_1
X_4512_ net1 VGND VPWR net38 u_usb_cdc.rstn_sq\[1\] clknet_leaf_19_clk_regs sg13g2_dfrbpq_1
Xhold104 _0208_ VPWR VGND net147 sg13g2_dlygate4sd3_1
XFILLER_8_693 VPWR VGND sg13g2_fill_1
Xhold126 _0100_ VPWR VGND net169 sg13g2_dlygate4sd3_1
Xhold115 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[32\] VPWR VGND
+ net158 sg13g2_dlygate4sd3_1
Xhold137 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[34\] VPWR
+ VGND net180 sg13g2_dlygate4sd3_1
Xhold148 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[67\] VPWR
+ VGND net191 sg13g2_dlygate4sd3_1
Xhold159 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[7\] VPWR VGND
+ net202 sg13g2_dlygate4sd3_1
X_4443_ net725 VGND VPWR net367 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[1\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_2
Xfanout606 net607 net606 VPWR VGND sg13g2_buf_1
X_4374_ net657 VGND VPWR _0302_ u_usb_cdc.bulk_out_nak[0] clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
X_3325_ VGND VPWR _1283_ _1323_ _0246_ net446 sg13g2_a21oi_1
Xfanout639 _0567_ net639 VPWR VGND sg13g2_buf_8
Xfanout617 _1284_ net617 VPWR VGND sg13g2_buf_8
Xfanout628 _1371_ net628 VPWR VGND sg13g2_buf_8
X_3256_ _1253_ _1258_ _1261_ _1262_ VPWR VGND sg13g2_nor3_1
X_2207_ net745 _0438_ _0439_ VPWR VGND sg13g2_and2_1
X_3187_ _1219_ VPWR _0212_ VGND net712 _1170_ sg13g2_o21ai_1
X_2138_ VPWR _1994_ net383 VGND sg13g2_inv_1
X_2069_ VPWR _1926_ u_usb_cdc.u_ctrl_endp.req_q\[2\] VGND sg13g2_inv_1
XFILLER_22_486 VPWR VGND sg13g2_fill_1
XFILLER_6_619 VPWR VGND sg13g2_decap_8
XFILLER_2_803 VPWR VGND sg13g2_decap_8
Xhold660 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] VPWR VGND net979 sg13g2_dlygate4sd3_1
Xhold671 _0051_ VPWR VGND net990 sg13g2_dlygate4sd3_1
Xhold693 u_usb_cdc.sie_out_data\[7\] VPWR VGND net1012 sg13g2_dlygate4sd3_1
XFILLER_1_346 VPWR VGND sg13g2_decap_8
Xhold682 u_usb_cdc.u_ctrl_endp.req_q\[9\] VPWR VGND net1001 sg13g2_dlygate4sd3_1
XFILLER_40_1013 VPWR VGND sg13g2_decap_8
XFILLER_40_1024 VPWR VGND sg13g2_fill_1
XFILLER_45_534 VPWR VGND sg13g2_fill_2
XFILLER_27_84 VPWR VGND sg13g2_fill_1
XFILLER_9_468 VPWR VGND sg13g2_fill_1
XFILLER_5_663 VPWR VGND sg13g2_decap_4
X_3110_ _1173_ net115 _1151_ VPWR VGND sg13g2_nand2_1
XFILLER_1_891 VPWR VGND sg13g2_decap_8
X_4090_ _1906_ VPWR _1907_ VGND net749 net551 sg13g2_o21ai_1
XFILLER_49_884 VPWR VGND sg13g2_decap_8
X_3041_ _1028_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\] _1031_
+ _1130_ VPWR VGND sg13g2_mux2_1
XFILLER_36_545 VPWR VGND sg13g2_fill_1
XFILLER_36_534 VPWR VGND sg13g2_decap_8
X_3943_ VGND VPWR _1796_ _1798_ _1799_ net707 sg13g2_a21oi_1
XFILLER_32_784 VPWR VGND sg13g2_fill_1
X_3874_ VGND VPWR net741 net361 _0370_ _1748_ sg13g2_a21oi_1
X_2825_ _0999_ u_usb_cdc.u_ctrl_endp.endp_q\[1\] u_usb_cdc.u_ctrl_endp.in_endp_q VPWR
+ VGND sg13g2_nand2_1
XFILLER_20_968 VPWR VGND sg13g2_fill_1
XFILLER_20_979 VPWR VGND sg13g2_decap_4
X_2756_ VGND VPWR net708 _0941_ _0047_ _0940_ sg13g2_a21oi_1
X_2687_ _1952_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[7\] _1949_ _0888_ VPWR VGND
+ _0887_ sg13g2_nand4_1
X_4426_ net684 VGND VPWR _0354_ u_usb_cdc.sie_out_data\[7\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_4357_ net686 VGND VPWR net954 u_usb_cdc.u_ctrl_endp.rec_q\[1\] clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_48_28 VPWR VGND sg13g2_decap_8
X_4288_ net673 VGND VPWR net417 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[50\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_3308_ VGND VPWR _1308_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[18\]
+ net823 sg13g2_or2_1
XFILLER_24_1019 VPWR VGND sg13g2_decap_8
X_3239_ _1247_ net166 _1156_ VPWR VGND sg13g2_nand2_1
XFILLER_27_567 VPWR VGND sg13g2_fill_1
XFILLER_27_556 VPWR VGND sg13g2_decap_8
XFILLER_42_537 VPWR VGND sg13g2_fill_2
XFILLER_11_968 VPWR VGND sg13g2_fill_1
Xhold490 _1812_ VPWR VGND net533 sg13g2_dlygate4sd3_1
XFILLER_49_125 VPWR VGND sg13g2_fill_2
XFILLER_18_512 VPWR VGND sg13g2_fill_2
XFILLER_46_876 VPWR VGND sg13g2_decap_8
XFILLER_18_578 VPWR VGND sg13g2_decap_4
XFILLER_18_589 VPWR VGND sg13g2_fill_2
XFILLER_14_784 VPWR VGND sg13g2_decap_8
X_3590_ _0338_ net580 _1496_ net584 _1953_ VPWR VGND sg13g2_a22oi_1
XFILLER_10_990 VPWR VGND sg13g2_decap_8
X_2610_ _0828_ net968 net591 VPWR VGND sg13g2_nand2_1
X_2541_ net721 net757 _0768_ VPWR VGND sg13g2_nor2_1
XFILLER_6_972 VPWR VGND sg13g2_decap_8
X_2472_ _0700_ _0637_ net623 VPWR VGND sg13g2_nand2_1
X_4211_ net666 VGND VPWR net518 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[57\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_4142_ net702 VGND VPWR net369 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_2
X_4073_ _1895_ net350 net389 VPWR VGND sg13g2_xnor2_1
X_3024_ _1120_ VPWR _0148_ VGND _1083_ _1098_ sg13g2_o21ai_1
XFILLER_49_681 VPWR VGND sg13g2_decap_8
X_3926_ _1746_ VPWR _1787_ VGND net352 _1783_ sg13g2_o21ai_1
XFILLER_32_581 VPWR VGND sg13g2_fill_1
X_3857_ _1735_ VPWR _0366_ VGND _1950_ net595 sg13g2_o21ai_1
X_2808_ _0984_ _0983_ u_usb_cdc.u_sie.in_toggle_q\[2\] _0514_ u_usb_cdc.u_sie.in_toggle_q\[0\]
+ VPWR VGND sg13g2_a22oi_1
X_3788_ _1687_ _1568_ u_usb_cdc.u_ctrl_endp.req_q\[2\] _1512_ _0660_ VPWR VGND sg13g2_a22oi_1
X_2739_ _0929_ net866 _0807_ VPWR VGND sg13g2_nand2_1
X_4409_ net696 VGND VPWR _0337_ u_usb_cdc.u_sie.crc16_q\[14\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_8_1013 VPWR VGND sg13g2_decap_8
X_4512__38 VPWR VGND net38 sg13g2_tiehi
XFILLER_28_810 VPWR VGND sg13g2_fill_2
XFILLER_42_312 VPWR VGND sg13g2_decap_8
XFILLER_15_537 VPWR VGND sg13g2_fill_2
XFILLER_42_378 VPWR VGND sg13g2_fill_1
XFILLER_10_253 VPWR VGND sg13g2_fill_2
XFILLER_11_765 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_8_clk_regs clknet_3_3__leaf_clk_regs clknet_leaf_8_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_40_40 VPWR VGND sg13g2_fill_2
XFILLER_3_975 VPWR VGND sg13g2_decap_8
XFILLER_49_82 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_fill_2
XFILLER_19_865 VPWR VGND sg13g2_fill_1
XFILLER_46_662 VPWR VGND sg13g2_decap_8
XFILLER_19_887 VPWR VGND sg13g2_decap_4
XFILLER_14_1007 VPWR VGND sg13g2_decap_8
X_3711_ _1613_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[68\] net628
+ VPWR VGND sg13g2_nand2_1
X_3642_ _1546_ VPWR _1547_ VGND _1441_ _1506_ sg13g2_o21ai_1
X_3573_ _0323_ net580 _1494_ net584 _1962_ VPWR VGND sg13g2_a22oi_1
X_2524_ u_usb_cdc.u_ctrl_endp.req_q\[2\] u_usb_cdc.u_ctrl_endp.req_q\[8\] _0751_ VPWR
+ VGND sg13g2_nor2_2
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_2455_ net787 _0669_ _0685_ VPWR VGND sg13g2_nor2_2
Xhold19 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[40\] VPWR VGND
+ net62 sg13g2_dlygate4sd3_1
X_2386_ _0611_ _0616_ _0617_ VPWR VGND sg13g2_nor2_2
X_4125_ net698 VGND VPWR _0026_ u_usb_cdc.u_sie.phy_state_q\[7\] clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_1
X_4056_ net308 _1842_ _1883_ VPWR VGND sg13g2_nor2_1
XFILLER_45_29 VPWR VGND sg13g2_fill_2
X_3007_ _1115_ net242 _1108_ VPWR VGND sg13g2_nand2_1
XFILLER_33_890 VPWR VGND sg13g2_fill_2
X_3909_ _1774_ net714 net340 VPWR VGND sg13g2_nand2_1
XFILLER_0_923 VPWR VGND sg13g2_decap_8
XFILLER_48_927 VPWR VGND sg13g2_decap_8
XFILLER_27_150 VPWR VGND sg13g2_fill_2
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_16_857 VPWR VGND sg13g2_fill_2
XFILLER_35_40 VPWR VGND sg13g2_decap_4
XFILLER_43_621 VPWR VGND sg13g2_decap_4
XFILLER_31_849 VPWR VGND sg13g2_fill_1
X_2240_ _0472_ u_usb_cdc.u_sie.data_q\[5\] _0458_ VPWR VGND sg13g2_xnor2_1
X_2171_ _0059_ _0058_ _0060_ _2027_ VPWR VGND sg13g2_nand3_1
XFILLER_20_1011 VPWR VGND sg13g2_decap_8
XFILLER_47_971 VPWR VGND sg13g2_decap_8
XFILLER_15_890 VPWR VGND sg13g2_fill_2
X_3625_ _1531_ _1528_ _1530_ VPWR VGND sg13g2_nand2_1
X_3556_ _1482_ net327 net598 VPWR VGND sg13g2_nand2_1
X_2507_ net880 net953 net794 _0734_ VPWR VGND sg13g2_nor3_1
X_3487_ _0619_ VPWR _1437_ VGND _0621_ _1436_ sg13g2_o21ai_1
XFILLER_5_1005 VPWR VGND sg13g2_decap_8
X_2438_ net791 net790 _0668_ VPWR VGND sg13g2_nor2_2
X_2369_ _0600_ net751 net840 VPWR VGND sg13g2_nand2_2
X_4108_ net687 VGND VPWR net858 u_usb_cdc.u_sie.in_toggle_q\[1\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_4039_ VPWR VGND _1868_ _1834_ _1823_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] _1869_
+ _0433_ sg13g2_a221oi_1
XFILLER_24_120 VPWR VGND sg13g2_fill_2
XFILLER_25_632 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_fill_1
XFILLER_25_665 VPWR VGND sg13g2_fill_1
XFILLER_9_809 VPWR VGND sg13g2_decap_4
XFILLER_21_893 VPWR VGND sg13g2_fill_2
XFILLER_0_720 VPWR VGND sg13g2_decap_8
XFILLER_0_797 VPWR VGND sg13g2_decap_8
XFILLER_48_724 VPWR VGND sg13g2_decap_8
XFILLER_44_963 VPWR VGND sg13g2_decap_8
Xhold308 _0422_ VPWR VGND net351 sg13g2_dlygate4sd3_1
X_3410_ VGND VPWR net724 net578 _0263_ _1391_ sg13g2_a21oi_1
X_4390_ net698 VGND VPWR net157 u_usb_cdc.u_sie.delay_cnt_q\[2\] clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_1
Xhold319 _0370_ VPWR VGND net362 sg13g2_dlygate4sd3_1
X_3341_ _1337_ VPWR _1338_ VGND _1288_ _1334_ sg13g2_o21ai_1
X_3272_ _1276_ _0604_ _1274_ net940 net755 VPWR VGND sg13g2_a22oi_1
X_2223_ _0455_ _0451_ _0454_ VPWR VGND sg13g2_nand2_1
X_2154_ VPWR _2010_ net23 VGND sg13g2_inv_1
X_2085_ VPWR _1942_ net1001 VGND sg13g2_inv_1
XFILLER_34_484 VPWR VGND sg13g2_decap_8
X_2987_ _1104_ VPWR _0127_ VGND _1052_ net610 sg13g2_o21ai_1
X_3608_ net788 net779 _0539_ _1514_ VPWR VGND sg13g2_nor3_2
XFILLER_1_539 VPWR VGND sg13g2_decap_8
X_3539_ _1470_ net955 _1466_ _0313_ VPWR VGND sg13g2_mux2_1
XFILLER_27_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_22_clk_regs clknet_3_6__leaf_clk_regs clknet_leaf_22_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_45_705 VPWR VGND sg13g2_decap_8
XFILLER_44_237 VPWR VGND sg13g2_fill_2
XFILLER_45_738 VPWR VGND sg13g2_decap_8
XFILLER_26_974 VPWR VGND sg13g2_decap_8
XFILLER_41_922 VPWR VGND sg13g2_fill_1
XFILLER_25_484 VPWR VGND sg13g2_fill_1
XFILLER_41_977 VPWR VGND sg13g2_decap_8
XFILLER_21_690 VPWR VGND sg13g2_fill_1
XFILLER_0_561 VPWR VGND sg13g2_decap_8
XFILLER_48_565 VPWR VGND sg13g2_decap_8
XFILLER_48_598 VPWR VGND sg13g2_decap_8
XFILLER_44_760 VPWR VGND sg13g2_decap_8
XFILLER_32_911 VPWR VGND sg13g2_decap_8
X_2910_ _1057_ net105 _1037_ VPWR VGND sg13g2_nand2_1
X_3890_ _1760_ net348 net387 _1754_ VPWR VGND sg13g2_and3_2
X_2841_ _1013_ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] net625 net747 _1909_ VPWR VGND
+ sg13g2_a22oi_1
X_2772_ net840 net839 _0950_ VPWR VGND sg13g2_nor2_1
XFILLER_8_661 VPWR VGND sg13g2_decap_4
X_4511_ net1 VGND VPWR net45 u_usb_cdc.rstn clknet_leaf_19_clk_regs sg13g2_dfrbpq_1
Xhold105 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[63\] VPWR
+ VGND net148 sg13g2_dlygate4sd3_1
Xhold116 _0115_ VPWR VGND net159 sg13g2_dlygate4sd3_1
X_4442_ net725 VGND VPWR net362 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[0\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_2
Xhold138 _0201_ VPWR VGND net181 sg13g2_dlygate4sd3_1
Xhold149 _0234_ VPWR VGND net192 sg13g2_dlygate4sd3_1
Xhold127 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[71\] VPWR
+ VGND net170 sg13g2_dlygate4sd3_1
X_4373_ net692 VGND VPWR net563 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] clknet_leaf_23_clk_regs
+ sg13g2_dfrbpq_2
X_3324_ _1323_ _1322_ _1983_ net629 net191 VPWR VGND sg13g2_a22oi_1
Xfanout629 _1294_ net629 VPWR VGND sg13g2_buf_8
Xfanout607 _1195_ net607 VPWR VGND sg13g2_buf_8
Xfanout618 net621 net618 VPWR VGND sg13g2_buf_8
X_3255_ _1259_ net820 _1261_ VPWR VGND sg13g2_xor2_1
X_2206_ _0438_ _0436_ _0435_ VPWR VGND sg13g2_nand2b_1
X_3186_ _1219_ net162 _1213_ VPWR VGND sg13g2_nand2_1
X_2137_ VPWR _1993_ net991 VGND sg13g2_inv_1
XFILLER_27_749 VPWR VGND sg13g2_decap_8
XFILLER_26_248 VPWR VGND sg13g2_fill_1
X_2068_ _1925_ net790 VPWR VGND sg13g2_inv_2
XFILLER_35_782 VPWR VGND sg13g2_fill_1
XFILLER_23_999 VPWR VGND sg13g2_decap_8
XFILLER_10_649 VPWR VGND sg13g2_fill_2
XFILLER_1_325 VPWR VGND sg13g2_decap_8
Xhold650 u_usb_cdc.u_ctrl_endp.state_q\[3\] VPWR VGND net969 sg13g2_dlygate4sd3_1
Xhold672 u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] VPWR VGND net991 sg13g2_dlygate4sd3_1
Xhold661 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\] VPWR VGND
+ net980 sg13g2_dlygate4sd3_1
XFILLER_2_859 VPWR VGND sg13g2_fill_1
Xhold694 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ VPWR VGND net1013 sg13g2_dlygate4sd3_1
Xhold683 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ VPWR VGND net1002 sg13g2_dlygate4sd3_1
XFILLER_27_63 VPWR VGND sg13g2_decap_8
XFILLER_45_513 VPWR VGND sg13g2_fill_1
XFILLER_45_557 VPWR VGND sg13g2_fill_1
XFILLER_14_933 VPWR VGND sg13g2_fill_1
XFILLER_43_40 VPWR VGND sg13g2_decap_8
XFILLER_40_262 VPWR VGND sg13g2_fill_2
XFILLER_9_458 VPWR VGND sg13g2_fill_1
XFILLER_5_686 VPWR VGND sg13g2_fill_1
XFILLER_49_863 VPWR VGND sg13g2_decap_8
X_3040_ net859 _1129_ _1128_ _0155_ VPWR VGND sg13g2_mux2_1
XFILLER_48_395 VPWR VGND sg13g2_decap_8
X_3942_ _1798_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] net423 VPWR VGND sg13g2_nand2_1
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
XFILLER_32_763 VPWR VGND sg13g2_fill_2
X_3873_ net361 net615 _1748_ VPWR VGND sg13g2_nor2_1
X_2824_ _0998_ _0997_ net378 _0992_ _0983_ VPWR VGND sg13g2_a22oi_1
XFILLER_9_981 VPWR VGND sg13g2_decap_8
X_2755_ _0941_ net567 net53 VPWR VGND sg13g2_nand2b_1
X_2686_ _0887_ _2036_ _2046_ _0886_ VPWR VGND sg13g2_and3_1
X_4425_ net684 VGND VPWR _0353_ u_usb_cdc.sie_out_data\[6\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_2
X_4356_ net686 VGND VPWR _0284_ u_usb_cdc.u_ctrl_endp.rec_q\[0\] clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_2
X_3307_ _1306_ VPWR _1307_ VGND net822 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[2\]
+ sg13g2_o21ai_1
X_4287_ net675 VGND VPWR net344 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[49\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
X_3238_ _1246_ VPWR _0236_ VGND _1155_ _1188_ sg13g2_o21ai_1
X_3169_ _1210_ net189 net608 VPWR VGND sg13g2_nand2_1
XFILLER_23_730 VPWR VGND sg13g2_fill_1
XFILLER_22_240 VPWR VGND sg13g2_fill_1
XFILLER_2_667 VPWR VGND sg13g2_decap_8
Xhold480 _0001_ VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold491 _0399_ VPWR VGND net534 sg13g2_dlygate4sd3_1
XFILLER_49_104 VPWR VGND sg13g2_decap_8
XFILLER_45_321 VPWR VGND sg13g2_fill_2
XFILLER_46_855 VPWR VGND sg13g2_decap_8
XFILLER_18_546 VPWR VGND sg13g2_fill_1
XFILLER_10_980 VPWR VGND sg13g2_fill_1
X_2540_ _0767_ _1936_ u_usb_cdc.u_ctrl_endp.rec_q\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_6_951 VPWR VGND sg13g2_decap_8
X_2471_ _0646_ _0662_ _1925_ _0699_ VPWR VGND net622 sg13g2_nand4_1
XFILLER_5_494 VPWR VGND sg13g2_decap_8
X_4210_ net667 VGND VPWR net508 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[56\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_4141_ net703 VGND VPWR _0036_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
X_4072_ _1894_ net389 net718 VPWR VGND sg13g2_nand2_1
XFILLER_23_1020 VPWR VGND sg13g2_decap_8
XFILLER_49_660 VPWR VGND sg13g2_decap_8
X_3023_ _1120_ net200 _1118_ VPWR VGND sg13g2_nand2_1
XFILLER_24_527 VPWR VGND sg13g2_fill_2
XFILLER_24_538 VPWR VGND sg13g2_decap_4
XFILLER_32_560 VPWR VGND sg13g2_fill_1
X_3925_ net352 _1783_ _1786_ VPWR VGND sg13g2_and2_1
X_3856_ _0899_ _1729_ net338 _1735_ VPWR VGND sg13g2_nand3_1
X_2807_ net768 u_usb_cdc.endp\[1\] _0983_ VPWR VGND sg13g2_nor2b_1
XFILLER_30_1024 VPWR VGND sg13g2_decap_4
X_3787_ VPWR _1686_ _1685_ VGND sg13g2_inv_1
X_2738_ VPWR _0038_ net925 VGND sg13g2_inv_1
X_4408_ net695 VGND VPWR net540 u_usb_cdc.u_sie.crc16_q\[13\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
X_2669_ net843 VPWR _0875_ VGND net598 _0874_ sg13g2_o21ai_1
X_4339_ net685 VGND VPWR _0267_ u_usb_cdc.u_ctrl_endp.in_endp_q clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_28_800 VPWR VGND sg13g2_fill_1
XFILLER_10_243 VPWR VGND sg13g2_fill_1
XFILLER_10_221 VPWR VGND sg13g2_fill_2
XFILLER_7_726 VPWR VGND sg13g2_decap_4
XFILLER_2_420 VPWR VGND sg13g2_fill_2
XFILLER_3_954 VPWR VGND sg13g2_decap_8
XFILLER_2_453 VPWR VGND sg13g2_decap_4
XFILLER_49_61 VPWR VGND sg13g2_decap_8
XFILLER_38_619 VPWR VGND sg13g2_fill_2
XFILLER_1_35 VPWR VGND sg13g2_decap_8
Xfanout790 net1052 net790 VPWR VGND sg13g2_buf_8
X_3710_ _1612_ VPWR _0342_ VGND _1610_ _1611_ sg13g2_o21ai_1
X_3641_ VGND VPWR _0533_ _1501_ _1546_ _1452_ sg13g2_a21oi_1
X_3572_ _1494_ _0497_ _0501_ VPWR VGND sg13g2_xnor2_1
X_2523_ u_usb_cdc.u_ctrl_endp.req_q\[1\] _0748_ _0749_ _0750_ VPWR VGND sg13g2_nor3_1
X_2454_ net759 net758 _0683_ _0684_ VPWR VGND sg13g2_nor3_1
X_2385_ _0614_ VPWR _0616_ VGND _0594_ _0606_ sg13g2_o21ai_1
X_4124_ net695 VGND VPWR net142 u_usb_cdc.u_sie.phy_state_q\[6\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_29_608 VPWR VGND sg13g2_decap_4
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_2
X_4055_ VPWR _0417_ net460 VGND sg13g2_inv_1
X_3006_ _1114_ VPWR _0136_ VGND _1072_ net611 sg13g2_o21ai_1
XFILLER_25_858 VPWR VGND sg13g2_fill_2
XFILLER_36_195 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_47_clk_regs clknet_3_1__leaf_clk_regs clknet_leaf_47_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3908_ _1771_ VPWR _0379_ VGND _1772_ _1773_ sg13g2_o21ai_1
X_3839_ _0359_ _1721_ _1724_ VPWR VGND sg13g2_nand2_1
XFILLER_3_206 VPWR VGND sg13g2_fill_1
XFILLER_0_902 VPWR VGND sg13g2_decap_8
XFILLER_48_906 VPWR VGND sg13g2_decap_8
XFILLER_0_979 VPWR VGND sg13g2_decap_8
XFILLER_19_20 VPWR VGND sg13g2_fill_1
XFILLER_31_817 VPWR VGND sg13g2_fill_1
XFILLER_3_773 VPWR VGND sg13g2_fill_1
X_2170_ _2026_ net1009 _0059_ _0058_ VPWR VGND sg13g2_and3_2
XFILLER_47_950 VPWR VGND sg13g2_decap_8
X_3624_ VGND VPWR net800 _1529_ _1530_ _1923_ sg13g2_a21oi_1
X_3555_ _0318_ _1481_ _1930_ _1475_ net746 VPWR VGND sg13g2_a22oi_1
X_2506_ _0709_ VPWR _0733_ VGND _1938_ _0722_ sg13g2_o21ai_1
X_3486_ net849 _1435_ _1436_ VPWR VGND sg13g2_nor2_1
X_2437_ net590 _0621_ _0666_ _0667_ VPWR VGND sg13g2_nor3_1
X_2368_ _0599_ net750 net752 VPWR VGND sg13g2_nand2b_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_4107_ net688 VGND VPWR net407 u_usb_cdc.u_sie.in_toggle_q\[0\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
X_2299_ _0524_ _0528_ _0529_ _0531_ VPWR VGND sg13g2_nor3_1
X_4038_ _1868_ _1866_ _1867_ VPWR VGND sg13g2_nand2_1
XFILLER_25_600 VPWR VGND sg13g2_fill_1
XFILLER_40_614 VPWR VGND sg13g2_fill_1
XFILLER_12_349 VPWR VGND sg13g2_decap_4
XFILLER_21_32 VPWR VGND sg13g2_decap_8
XFILLER_4_559 VPWR VGND sg13g2_fill_1
XFILLER_48_703 VPWR VGND sg13g2_decap_8
XFILLER_0_776 VPWR VGND sg13g2_decap_8
XFILLER_46_40 VPWR VGND sg13g2_decap_8
XFILLER_44_942 VPWR VGND sg13g2_decap_8
XFILLER_29_994 VPWR VGND sg13g2_decap_8
XFILLER_16_644 VPWR VGND sg13g2_fill_2
XFILLER_16_688 VPWR VGND sg13g2_decap_4
XFILLER_31_603 VPWR VGND sg13g2_fill_2
XFILLER_43_496 VPWR VGND sg13g2_fill_1
XFILLER_8_810 VPWR VGND sg13g2_fill_1
XFILLER_7_34 VPWR VGND sg13g2_fill_1
XFILLER_7_67 VPWR VGND sg13g2_fill_1
XFILLER_8_876 VPWR VGND sg13g2_fill_1
Xhold309 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[14\] VPWR VGND net352 sg13g2_dlygate4sd3_1
X_3340_ _1337_ _1335_ _1336_ _1332_ net812 VPWR VGND sg13g2_a22oi_1
X_3271_ _1275_ _0714_ _1256_ VPWR VGND sg13g2_nand2_1
XFILLER_30_4 VPWR VGND sg13g2_decap_8
X_2222_ _1934_ net1028 _0454_ VPWR VGND sg13g2_nor2_1
X_2153_ VPWR _2009_ net259 VGND sg13g2_inv_1
XFILLER_16_2 VPWR VGND sg13g2_fill_1
X_2084_ VPWR _1941_ u_usb_cdc.u_ctrl_endp.req_q\[7\] VGND sg13g2_inv_1
XFILLER_35_997 VPWR VGND sg13g2_decap_8
XFILLER_22_625 VPWR VGND sg13g2_fill_1
X_2986_ _1104_ net90 _1096_ VPWR VGND sg13g2_nand2_1
X_3607_ _1513_ u_usb_cdc.u_ctrl_endp.req_q\[8\] net772 VPWR VGND sg13g2_nand2b_1
X_3538_ _1469_ VPWR _1470_ VGND net489 _1940_ sg13g2_o21ai_1
XFILLER_1_518 VPWR VGND sg13g2_decap_8
X_3469_ VGND VPWR net576 _1424_ _0289_ _1423_ sg13g2_a21oi_1
XFILLER_29_246 VPWR VGND sg13g2_fill_2
XFILLER_44_227 VPWR VGND sg13g2_fill_1
XFILLER_41_956 VPWR VGND sg13g2_decap_8
XFILLER_20_190 VPWR VGND sg13g2_fill_1
XFILLER_5_835 VPWR VGND sg13g2_fill_1
XFILLER_10_1011 VPWR VGND sg13g2_decap_8
XFILLER_0_540 VPWR VGND sg13g2_decap_8
XFILLER_48_544 VPWR VGND sg13g2_fill_2
XFILLER_17_964 VPWR VGND sg13g2_fill_1
X_2840_ VGND VPWR _1010_ _1011_ _1012_ _2022_ sg13g2_a21oi_1
XFILLER_43_282 VPWR VGND sg13g2_fill_2
XFILLER_32_989 VPWR VGND sg13g2_decap_8
X_2771_ _0949_ _0841_ _0947_ _0948_ VPWR VGND sg13g2_and3_1
XFILLER_8_651 VPWR VGND sg13g2_fill_2
X_4510_ net731 VGND VPWR _0040_ u_usb_cdc.clk_cnt_q\[1\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
X_4441_ net735 VGND VPWR _0369_ _0056_ clknet_leaf_26_clk_regs sg13g2_dfrbpq_2
Xhold117 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[30\] VPWR
+ VGND net160 sg13g2_dlygate4sd3_1
Xhold106 _0230_ VPWR VGND net149 sg13g2_dlygate4sd3_1
Xhold128 _0238_ VPWR VGND net171 sg13g2_dlygate4sd3_1
Xhold139 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[18\] VPWR VGND
+ net182 sg13g2_dlygate4sd3_1
X_4372_ net694 VGND VPWR _0300_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[5\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_1
Xfanout608 net609 net608 VPWR VGND sg13g2_buf_8
X_3323_ _1322_ _1319_ _1321_ _1317_ _1315_ VPWR VGND sg13g2_a22oi_1
Xfanout619 net621 net619 VPWR VGND sg13g2_buf_8
X_3254_ VPWR _1260_ _1259_ VGND sg13g2_inv_1
X_2205_ VPWR _0437_ _0436_ VGND sg13g2_inv_1
X_3185_ _1218_ VPWR _0211_ VGND net712 _1168_ sg13g2_o21ai_1
X_2136_ VPWR _1992_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[15\]
+ VGND sg13g2_inv_1
X_2067_ _1924_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\]
+ VPWR VGND sg13g2_inv_2
XFILLER_10_606 VPWR VGND sg13g2_decap_8
X_2969_ _1093_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net636 VPWR VGND sg13g2_nand2_1
XFILLER_1_304 VPWR VGND sg13g2_fill_1
Xhold640 u_usb_cdc.u_ctrl_endp.state_q\[1\] VPWR VGND net959 sg13g2_dlygate4sd3_1
Xhold651 _0013_ VPWR VGND net970 sg13g2_dlygate4sd3_1
Xhold662 _0262_ VPWR VGND net981 sg13g2_dlygate4sd3_1
Xhold684 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[0\] VPWR VGND
+ net1003 sg13g2_dlygate4sd3_1
Xhold673 u_usb_cdc.u_sie.data_q\[6\] VPWR VGND net992 sg13g2_dlygate4sd3_1
Xhold695 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[1\] VPWR VGND
+ net1014 sg13g2_dlygate4sd3_1
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_14_901 VPWR VGND sg13g2_decap_8
XFILLER_49_842 VPWR VGND sg13g2_decap_8
X_3941_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\] u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\]
+ _1797_ VPWR VGND sg13g2_and2_1
XFILLER_16_282 VPWR VGND sg13g2_fill_2
XFILLER_17_1006 VPWR VGND sg13g2_decap_8
XFILLER_32_753 VPWR VGND sg13g2_decap_4
X_3872_ _1747_ net744 VPWR VGND _1745_ sg13g2_nand2b_2
X_2823_ _0997_ _0987_ _0996_ VPWR VGND sg13g2_nand2_1
X_2754_ net53 _0940_ _0046_ VPWR VGND sg13g2_nor2_1
X_2685_ _0056_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] net312 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\]
+ _0886_ VPWR VGND sg13g2_nor4_1
X_4424_ net684 VGND VPWR _0352_ u_usb_cdc.sie_out_data\[5\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_2
X_4355_ net690 VGND VPWR _0283_ u_usb_cdc.u_ctrl_endp.dev_state_q\[1\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_3306_ _1306_ net822 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[10\]
+ VPWR VGND sg13g2_nand2b_1
X_4286_ net675 VGND VPWR net318 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[48\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
X_3237_ _1246_ net226 _1156_ VPWR VGND sg13g2_nand2_1
X_3168_ _1209_ VPWR _0203_ VGND _1186_ net608 sg13g2_o21ai_1
X_2119_ VPWR _1976_ net274 VGND sg13g2_inv_1
X_3099_ net830 _1159_ net760 _1166_ VPWR VGND sg13g2_nand3_1
XFILLER_11_915 VPWR VGND sg13g2_decap_8
XFILLER_11_926 VPWR VGND sg13g2_fill_1
XFILLER_13_55 VPWR VGND sg13g2_fill_2
Xhold481 u_usb_cdc.u_sie.phy_state_q\[2\] VPWR VGND net524 sg13g2_dlygate4sd3_1
XFILLER_2_646 VPWR VGND sg13g2_fill_1
Xhold470 u_usb_cdc.u_ctrl_endp.req_q\[5\] VPWR VGND net513 sg13g2_dlygate4sd3_1
Xhold492 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[28\] VPWR VGND
+ net535 sg13g2_dlygate4sd3_1
XFILLER_49_127 VPWR VGND sg13g2_fill_1
XFILLER_46_834 VPWR VGND sg13g2_decap_8
XFILLER_18_514 VPWR VGND sg13g2_fill_1
XFILLER_38_96 VPWR VGND sg13g2_fill_2
XFILLER_45_300 VPWR VGND sg13g2_decap_4
XFILLER_45_377 VPWR VGND sg13g2_fill_1
XFILLER_41_561 VPWR VGND sg13g2_fill_1
X_2470_ _0698_ net723 _0692_ VPWR VGND sg13g2_nand2_1
XFILLER_5_473 VPWR VGND sg13g2_decap_8
X_4140_ net702 VGND VPWR _0066_ _0053_ clknet_leaf_37_clk_regs sg13g2_dfrbpq_2
X_4071_ _1893_ VPWR _0422_ VGND net350 _1892_ sg13g2_o21ai_1
X_3022_ _1119_ VPWR _0147_ VGND _1081_ _1098_ sg13g2_o21ai_1
XFILLER_48_160 VPWR VGND sg13g2_fill_2
XFILLER_17_580 VPWR VGND sg13g2_decap_8
X_3924_ _1785_ net714 net352 VPWR VGND sg13g2_nand2_1
X_3855_ _1734_ VPWR _0365_ VGND _1951_ net595 sg13g2_o21ai_1
X_2806_ _0982_ u_usb_cdc.u_sie.in_toggle_q\[1\] _0566_ VPWR VGND sg13g2_nand2_1
XFILLER_30_1003 VPWR VGND sg13g2_decap_8
X_3786_ _1685_ _1683_ _1684_ net628 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[71\]
+ VPWR VGND sg13g2_a22oi_1
X_2737_ _0928_ _0924_ net924 _0923_ net835 VPWR VGND sg13g2_a22oi_1
X_2668_ net753 _0556_ _0564_ _0585_ _0874_ VPWR VGND sg13g2_nor4_1
X_4407_ net700 VGND VPWR net914 u_usb_cdc.u_sie.crc16_q\[12\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
X_2599_ u_usb_cdc.u_ctrl_endp.max_length_q\[4\] u_usb_cdc.u_ctrl_endp.max_length_q\[5\]
+ u_usb_cdc.u_ctrl_endp.max_length_q\[6\] _0818_ VPWR VGND sg13g2_nor3_1
X_4338_ net683 VGND VPWR _0266_ u_usb_cdc.u_ctrl_endp.endp_q\[3\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
X_4269_ net674 VGND VPWR net371 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[31\]
+ clknet_leaf_47_clk_regs sg13g2_dfrbpq_1
XFILLER_28_834 VPWR VGND sg13g2_fill_1
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_24_54 VPWR VGND sg13g2_decap_8
XFILLER_11_756 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_fill_1
XFILLER_40_97 VPWR VGND sg13g2_fill_2
XFILLER_49_40 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
Xfanout791 net793 net791 VPWR VGND sg13g2_buf_8
Xfanout780 net781 net780 VPWR VGND sg13g2_buf_8
XFILLER_1_58 VPWR VGND sg13g2_fill_1
XFILLER_46_697 VPWR VGND sg13g2_decap_8
X_3640_ _1543_ VPWR _1545_ VGND net781 _1544_ sg13g2_o21ai_1
X_3571_ net847 net921 net584 _1493_ VPWR VGND sg13g2_nor3_2
X_2522_ VGND VPWR _0749_ u_usb_cdc.u_ctrl_endp.req_q\[11\] u_usb_cdc.u_ctrl_endp.req_q\[4\]
+ sg13g2_or2_1
X_2453_ _0682_ VPWR _0683_ VGND net723 net721 sg13g2_o21ai_1
X_2384_ _0615_ _0612_ _0613_ VPWR VGND sg13g2_nand2_2
X_4123_ net688 VGND VPWR net302 u_usb_cdc.u_sie.phy_state_q\[5\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
X_4054_ _1882_ _1842_ _1881_ net642 net459 VPWR VGND sg13g2_a22oi_1
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
X_3005_ _1114_ net240 _1108_ VPWR VGND sg13g2_nand2_1
X_3907_ net615 VPWR _1773_ VGND net391 _1769_ sg13g2_o21ai_1
X_3838_ net745 _0437_ net840 _1724_ VPWR VGND _1723_ sg13g2_nand4_1
Xclkbuf_leaf_16_clk_regs clknet_3_2__leaf_clk_regs clknet_leaf_16_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3769_ _1661_ VPWR _1669_ VGND net795 _1668_ sg13g2_o21ai_1
XFILLER_0_958 VPWR VGND sg13g2_decap_8
XFILLER_19_119 VPWR VGND sg13g2_fill_2
XFILLER_28_620 VPWR VGND sg13g2_decap_8
XFILLER_43_645 VPWR VGND sg13g2_fill_2
XFILLER_24_892 VPWR VGND sg13g2_decap_4
XFILLER_24_881 VPWR VGND sg13g2_fill_2
XFILLER_19_631 VPWR VGND sg13g2_decap_8
XFILLER_34_601 VPWR VGND sg13g2_fill_1
XFILLER_46_483 VPWR VGND sg13g2_fill_1
XFILLER_34_667 VPWR VGND sg13g2_decap_8
XFILLER_30_840 VPWR VGND sg13g2_fill_1
X_3623_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[48\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[56\]
+ net807 _1529_ VPWR VGND sg13g2_mux2_1
X_3554_ u_usb_cdc.u_sie.delay_cnt_q\[0\] net745 u_usb_cdc.u_sie.delay_cnt_q\[1\] _1481_
+ VPWR VGND sg13g2_nand3_1
X_2505_ _0732_ _1938_ _0706_ VPWR VGND sg13g2_nand2_1
X_3485_ VGND VPWR _0549_ _0624_ _1435_ _1929_ sg13g2_a21oi_1
X_2436_ _0666_ net850 _0602_ VPWR VGND sg13g2_nand2_1
X_2367_ VPWR VGND _0597_ _0516_ _0596_ _0592_ _0598_ _0593_ sg13g2_a221oi_1
X_2298_ net790 u_usb_cdc.u_ctrl_endp.max_length_q\[1\] _0530_ VPWR VGND sg13g2_xor2_1
X_4106_ net689 VGND VPWR net56 u_usb_cdc.u_sie.out_toggle_q\[1\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_1
X_4037_ _1867_ u_usb_cdc.u_sie.data_q\[5\] net843 _1933_ u_usb_cdc.u_sie.phy_state_q\[11\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_38_995 VPWR VGND sg13g2_decap_8
XFILLER_25_689 VPWR VGND sg13g2_fill_2
XFILLER_24_199 VPWR VGND sg13g2_fill_1
XFILLER_43_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_755 VPWR VGND sg13g2_decap_8
XFILLER_48_759 VPWR VGND sg13g2_decap_8
XFILLER_29_973 VPWR VGND sg13g2_decap_8
XFILLER_44_921 VPWR VGND sg13g2_decap_8
XFILLER_44_998 VPWR VGND sg13g2_decap_8
X_3270_ _1273_ VPWR _1274_ VGND net770 net711 sg13g2_o21ai_1
X_2221_ net998 _0450_ _0452_ _0453_ VPWR VGND sg13g2_or3_1
XFILLER_23_4 VPWR VGND sg13g2_decap_8
X_2152_ VPWR _2008_ net296 VGND sg13g2_inv_1
X_2083_ _1940_ net851 VPWR VGND sg13g2_inv_2
XFILLER_35_976 VPWR VGND sg13g2_decap_8
XFILLER_22_637 VPWR VGND sg13g2_decap_8
XFILLER_21_147 VPWR VGND sg13g2_fill_2
X_2985_ _1103_ VPWR _0126_ VGND _1050_ net610 sg13g2_o21ai_1
X_3606_ net772 u_usb_cdc.u_ctrl_endp.req_q\[8\] _1512_ VPWR VGND sg13g2_nor2b_1
X_3537_ VGND VPWR net917 _1469_ _1468_ _1467_ sg13g2_a21oi_2
X_3468_ u_usb_cdc.sie_out_data\[1\] _1421_ _1424_ VPWR VGND sg13g2_nor2_1
X_2419_ _0649_ net743 _0648_ VPWR VGND sg13g2_nand2_1
X_3399_ _1369_ _1382_ _1383_ VPWR VGND sg13g2_nor2_1
XFILLER_26_921 VPWR VGND sg13g2_fill_2
XFILLER_26_910 VPWR VGND sg13g2_fill_2
XFILLER_41_935 VPWR VGND sg13g2_decap_8
XFILLER_13_626 VPWR VGND sg13g2_decap_4
XFILLER_16_99 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_31_clk_regs clknet_3_7__leaf_clk_regs clknet_leaf_31_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_5_858 VPWR VGND sg13g2_decap_8
XFILLER_5_869 VPWR VGND sg13g2_fill_1
XFILLER_0_596 VPWR VGND sg13g2_fill_2
XFILLER_48_523 VPWR VGND sg13g2_decap_8
XFILLER_32_968 VPWR VGND sg13g2_decap_8
X_2770_ _0450_ _0479_ net838 _0948_ VPWR VGND sg13g2_nand3_1
XFILLER_8_641 VPWR VGND sg13g2_fill_1
XFILLER_8_685 VPWR VGND sg13g2_fill_2
X_4440_ net730 VGND VPWR net964 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[7\] clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_2
Xhold107 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[55\] VPWR VGND
+ net150 sg13g2_dlygate4sd3_1
Xhold129 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[24\] VPWR
+ VGND net172 sg13g2_dlygate4sd3_1
Xhold118 _0197_ VPWR VGND net161 sg13g2_dlygate4sd3_1
X_4371_ net692 VGND VPWR _0299_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[4\] clknet_leaf_23_clk_regs
+ sg13g2_dfrbpq_1
X_3322_ VGND VPWR net816 _1320_ _1321_ _1982_ sg13g2_a21oi_1
Xfanout609 _1204_ net609 VPWR VGND sg13g2_buf_8
X_3253_ VGND VPWR net826 _1154_ _1259_ net831 sg13g2_a21oi_1
X_3184_ _1218_ net230 _1213_ VPWR VGND sg13g2_nand2_1
X_2204_ net751 net753 net465 _0436_ VPWR VGND sg13g2_nor3_2
XFILLER_39_534 VPWR VGND sg13g2_fill_1
X_2135_ VPWR _1991_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[46\]
+ VGND sg13g2_inv_1
X_2066_ net797 _1923_ VPWR VGND sg13g2_inv_4
XFILLER_35_773 VPWR VGND sg13g2_fill_2
XFILLER_23_968 VPWR VGND sg13g2_decap_8
XFILLER_33_1012 VPWR VGND sg13g2_decap_8
XFILLER_33_1023 VPWR VGND sg13g2_fill_2
X_2968_ _1092_ net196 _1079_ VPWR VGND sg13g2_nand2_1
X_2899_ _1050_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net645 VPWR VGND sg13g2_nand2_1
Xhold630 u_usb_cdc.u_ctrl_endp.state_q\[7\] VPWR VGND net949 sg13g2_dlygate4sd3_1
Xhold652 u_usb_cdc.endp\[3\] VPWR VGND net971 sg13g2_dlygate4sd3_1
XFILLER_2_839 VPWR VGND sg13g2_fill_2
Xhold641 _0011_ VPWR VGND net960 sg13g2_dlygate4sd3_1
Xhold663 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[3\] VPWR VGND net982 sg13g2_dlygate4sd3_1
Xhold674 u_usb_cdc.endp\[0\] VPWR VGND net993 sg13g2_dlygate4sd3_1
Xhold685 _0251_ VPWR VGND net1004 sg13g2_dlygate4sd3_1
Xhold696 _1377_ VPWR VGND net1015 sg13g2_dlygate4sd3_1
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_27_98 VPWR VGND sg13g2_fill_1
XFILLER_32_209 VPWR VGND sg13g2_fill_2
XFILLER_14_979 VPWR VGND sg13g2_fill_1
XFILLER_41_765 VPWR VGND sg13g2_decap_4
XFILLER_4_198 VPWR VGND sg13g2_fill_1
XFILLER_49_821 VPWR VGND sg13g2_decap_8
XFILLER_0_393 VPWR VGND sg13g2_decap_8
XFILLER_49_898 VPWR VGND sg13g2_decap_8
XFILLER_1_1010 VPWR VGND sg13g2_decap_8
X_3940_ _1796_ net707 net979 _0388_ VPWR VGND sg13g2_mux2_1
X_3871_ net713 _1745_ _1746_ VPWR VGND sg13g2_nor2_2
X_2822_ _2014_ _0983_ _0996_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_961 VPWR VGND sg13g2_fill_2
X_2753_ _0940_ _0938_ _0939_ VPWR VGND sg13g2_nand2_1
X_2684_ _0883_ VPWR _0885_ VGND _2035_ _0884_ sg13g2_o21ai_1
X_4423_ net684 VGND VPWR _0351_ u_usb_cdc.sie_out_data\[4\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_2
X_4354_ net690 VGND VPWR _0282_ _0055_ clknet_leaf_44_clk_regs sg13g2_dfrbpq_1
X_3305_ net821 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[34\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[42\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[50\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[58\] net816 _1305_
+ VPWR VGND sg13g2_mux4_1
X_4285_ net657 VGND VPWR net99 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[47\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
X_3236_ _1245_ VPWR _0235_ VGND _1155_ _1186_ sg13g2_o21ai_1
XFILLER_39_353 VPWR VGND sg13g2_decap_4
X_3167_ _1209_ net185 net608 VPWR VGND sg13g2_nand2_1
X_2118_ VPWR _1975_ net961 VGND sg13g2_inv_1
X_3098_ _1165_ net278 _1151_ VPWR VGND sg13g2_nand2_1
XFILLER_10_426 VPWR VGND sg13g2_decap_8
Xhold471 _0006_ VPWR VGND net514 sg13g2_dlygate4sd3_1
XFILLER_2_625 VPWR VGND sg13g2_fill_1
Xhold460 _0043_ VPWR VGND net503 sg13g2_dlygate4sd3_1
XFILLER_1_146 VPWR VGND sg13g2_fill_2
Xhold482 _0021_ VPWR VGND net525 sg13g2_dlygate4sd3_1
Xhold493 _0111_ VPWR VGND net536 sg13g2_dlygate4sd3_1
XFILLER_46_802 VPWR VGND sg13g2_decap_8
XFILLER_14_754 VPWR VGND sg13g2_fill_2
XFILLER_9_213 VPWR VGND sg13g2_fill_2
XFILLER_41_584 VPWR VGND sg13g2_fill_2
XFILLER_9_279 VPWR VGND sg13g2_fill_2
XFILLER_6_986 VPWR VGND sg13g2_decap_8
X_4070_ _1893_ net350 net718 VPWR VGND sg13g2_nand2_1
X_3021_ _1119_ net92 _1118_ VPWR VGND sg13g2_nand2_1
XFILLER_49_695 VPWR VGND sg13g2_decap_8
XFILLER_45_890 VPWR VGND sg13g2_decap_8
X_3923_ _1782_ VPWR _0383_ VGND _1783_ _1784_ sg13g2_o21ai_1
X_3854_ _0899_ _1729_ net310 _1734_ VPWR VGND sg13g2_nand3_1
X_2805_ net406 VPWR _0981_ VGND _0516_ _0980_ sg13g2_o21ai_1
X_3785_ VGND VPWR _1676_ _1678_ _1684_ net795 sg13g2_a21oi_1
X_2736_ _0927_ VPWR _0037_ VGND net368 _2025_ sg13g2_o21ai_1
X_2667_ _0873_ VPWR _0025_ VGND net141 _0844_ sg13g2_o21ai_1
X_4406_ net700 VGND VPWR net903 u_usb_cdc.u_sie.crc16_q\[11\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
X_2598_ VGND VPWR _0595_ _0617_ _0817_ net591 sg13g2_a21oi_1
X_4337_ net683 VGND VPWR net546 u_usb_cdc.u_ctrl_endp.endp_q\[2\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_8_1027 VPWR VGND sg13g2_fill_2
X_4268_ net656 VGND VPWR net161 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[30\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_3219_ _1237_ net303 net603 VPWR VGND sg13g2_nand2_1
XFILLER_28_857 VPWR VGND sg13g2_fill_2
X_4199_ net662 VGND VPWR net118 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[45\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
XFILLER_39_194 VPWR VGND sg13g2_fill_1
XFILLER_42_326 VPWR VGND sg13g2_fill_1
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_10_234 VPWR VGND sg13g2_fill_2
XFILLER_10_223 VPWR VGND sg13g2_fill_1
XFILLER_11_779 VPWR VGND sg13g2_fill_1
XFILLER_6_249 VPWR VGND sg13g2_fill_2
XFILLER_2_400 VPWR VGND sg13g2_decap_8
XFILLER_2_466 VPWR VGND sg13g2_decap_4
XFILLER_3_989 VPWR VGND sg13g2_decap_8
Xhold290 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[23\] VPWR
+ VGND net333 sg13g2_dlygate4sd3_1
Xfanout770 net771 net770 VPWR VGND sg13g2_buf_8
XFILLER_19_824 VPWR VGND sg13g2_fill_1
Xfanout792 net793 net792 VPWR VGND sg13g2_buf_1
Xfanout781 net782 net781 VPWR VGND sg13g2_buf_8
XFILLER_46_676 VPWR VGND sg13g2_decap_8
X_3570_ _1492_ net594 _1491_ VPWR VGND sg13g2_nand2_2
X_2521_ _0748_ _1941_ _0747_ VPWR VGND sg13g2_nand2_1
X_2452_ net760 net761 _0682_ VPWR VGND sg13g2_nor2_2
X_2383_ _0612_ _0613_ _0614_ VPWR VGND sg13g2_and2_1
X_4122_ net697 VGND VPWR _0023_ u_usb_cdc.u_sie.phy_state_q\[4\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_1
X_4053_ _1881_ _1832_ _1880_ net709 net835 VPWR VGND sg13g2_a22oi_1
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
X_3004_ _1113_ VPWR _0135_ VGND _1070_ net611 sg13g2_o21ai_1
XFILLER_49_492 VPWR VGND sg13g2_decap_8
XFILLER_25_849 VPWR VGND sg13g2_fill_2
X_3906_ net391 _1769_ _1772_ VPWR VGND sg13g2_and2_1
X_3837_ _0713_ VPWR _1723_ VGND _0506_ _1722_ sg13g2_o21ai_1
X_3768_ _1667_ VPWR _1668_ VGND net797 _1662_ sg13g2_o21ai_1
X_2719_ _0915_ VPWR _0032_ VGND _0881_ _0888_ sg13g2_o21ai_1
X_3699_ _1602_ u_usb_cdc.u_ctrl_endp.req_q\[8\] _0537_ VPWR VGND sg13g2_nand2_1
XFILLER_0_937 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_27_175 VPWR VGND sg13g2_fill_2
XFILLER_13_1010 VPWR VGND sg13g2_decap_8
XFILLER_7_547 VPWR VGND sg13g2_fill_2
XFILLER_3_731 VPWR VGND sg13g2_decap_8
XFILLER_3_742 VPWR VGND sg13g2_fill_2
XFILLER_47_985 VPWR VGND sg13g2_decap_8
XFILLER_18_142 VPWR VGND sg13g2_fill_1
XFILLER_19_665 VPWR VGND sg13g2_fill_2
XFILLER_20_1025 VPWR VGND sg13g2_decap_4
XFILLER_46_451 VPWR VGND sg13g2_fill_1
XFILLER_34_635 VPWR VGND sg13g2_fill_2
XFILLER_34_657 VPWR VGND sg13g2_fill_2
XFILLER_30_863 VPWR VGND sg13g2_fill_2
X_3622_ _1527_ VPWR _1528_ VGND net810 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[32\]
+ sg13g2_o21ai_1
X_3553_ net431 VPWR _0317_ VGND _1477_ _1480_ sg13g2_o21ai_1
X_2504_ _0731_ _0730_ _0725_ VPWR VGND sg13g2_nand2b_1
X_3484_ VGND VPWR net577 _1434_ _0294_ _1433_ sg13g2_a21oi_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_2435_ _0601_ net850 _0665_ VPWR VGND sg13g2_nor2b_2
X_4105_ net686 VGND VPWR net523 u_usb_cdc.u_ctrl_endp.req_q\[11\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_5_1019 VPWR VGND sg13g2_decap_8
X_2366_ VGND VPWR _1918_ u_usb_cdc.u_ctrl_endp.state_q\[3\] _0597_ u_usb_cdc.u_ctrl_endp.state_q\[2\]
+ sg13g2_a21oi_1
X_2297_ net775 u_usb_cdc.u_ctrl_endp.max_length_q\[5\] _0529_ VPWR VGND sg13g2_xor2_1
XFILLER_38_974 VPWR VGND sg13g2_decap_8
XFILLER_38_963 VPWR VGND sg13g2_fill_2
X_4036_ _1866_ _1965_ net837 _1958_ net846 VPWR VGND sg13g2_a22oi_1
XFILLER_36_1021 VPWR VGND sg13g2_decap_8
XFILLER_21_830 VPWR VGND sg13g2_fill_1
XFILLER_43_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_734 VPWR VGND sg13g2_decap_8
XFILLER_48_738 VPWR VGND sg13g2_decap_8
XFILLER_44_900 VPWR VGND sg13g2_decap_8
XFILLER_29_952 VPWR VGND sg13g2_decap_8
XFILLER_28_484 VPWR VGND sg13g2_fill_1
XFILLER_44_977 VPWR VGND sg13g2_decap_8
XFILLER_16_668 VPWR VGND sg13g2_fill_2
XFILLER_15_167 VPWR VGND sg13g2_fill_1
XFILLER_15_145 VPWR VGND sg13g2_fill_2
XFILLER_31_638 VPWR VGND sg13g2_decap_8
XFILLER_8_801 VPWR VGND sg13g2_decap_8
XFILLER_8_834 VPWR VGND sg13g2_fill_1
XFILLER_3_561 VPWR VGND sg13g2_decap_8
X_2220_ _0452_ u_usb_cdc.u_sie.pid_q\[3\] _0451_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_1_clk_regs clknet_3_0__leaf_clk_regs clknet_leaf_1_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2151_ VPWR _2007_ net368 VGND sg13g2_inv_1
X_2082_ net744 _1939_ VPWR VGND sg13g2_inv_4
XFILLER_47_782 VPWR VGND sg13g2_decap_8
XFILLER_35_911 VPWR VGND sg13g2_fill_1
XFILLER_19_484 VPWR VGND sg13g2_fill_2
XFILLER_34_498 VPWR VGND sg13g2_decap_8
X_2984_ _1103_ net59 _1096_ VPWR VGND sg13g2_nand2_1
XFILLER_30_671 VPWR VGND sg13g2_fill_1
X_3605_ VGND VPWR _0647_ _0669_ _1511_ _1452_ sg13g2_a21oi_1
X_3536_ net851 u_usb_cdc.u_ctrl_endp.addr_dd\[1\] u_usb_cdc.u_ctrl_endp.addr_dd\[0\]
+ u_usb_cdc.u_ctrl_endp.addr_dd\[3\] _1468_ VPWR VGND sg13g2_nor4_1
X_3467_ net926 net576 _1423_ VPWR VGND sg13g2_nor2_1
X_2418_ _0534_ _0645_ _0648_ VPWR VGND sg13g2_nor2_1
X_3398_ VGND VPWR _1133_ _1381_ _1382_ _1378_ sg13g2_a21oi_1
X_2349_ VGND VPWR _0518_ net987 _0581_ net596 sg13g2_a21oi_1
XFILLER_29_248 VPWR VGND sg13g2_fill_1
XFILLER_45_719 VPWR VGND sg13g2_decap_8
X_4019_ net626 _2026_ _1849_ _1850_ _1851_ VPWR VGND sg13g2_and4_1
XFILLER_41_903 VPWR VGND sg13g2_decap_8
XFILLER_16_78 VPWR VGND sg13g2_decap_4
XFILLER_26_988 VPWR VGND sg13g2_decap_8
XFILLER_9_609 VPWR VGND sg13g2_fill_1
XFILLER_21_671 VPWR VGND sg13g2_fill_2
XFILLER_5_815 VPWR VGND sg13g2_fill_2
XFILLER_4_347 VPWR VGND sg13g2_decap_4
XFILLER_4_369 VPWR VGND sg13g2_decap_4
XFILLER_0_575 VPWR VGND sg13g2_decap_8
XFILLER_48_513 VPWR VGND sg13g2_fill_1
XFILLER_48_557 VPWR VGND sg13g2_fill_2
XFILLER_32_925 VPWR VGND sg13g2_decap_8
XFILLER_44_774 VPWR VGND sg13g2_decap_8
XFILLER_32_958 VPWR VGND sg13g2_fill_1
XFILLER_12_671 VPWR VGND sg13g2_fill_2
Xhold108 _0138_ VPWR VGND net151 sg13g2_dlygate4sd3_1
Xhold119 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[45\] VPWR
+ VGND net162 sg13g2_dlygate4sd3_1
Xheichips25_usb_cdc_40 VPWR VGND uio_oe[4] sg13g2_tiehi
X_4370_ net694 VGND VPWR _0298_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[3\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_1
X_3321_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[51\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[59\]
+ net821 _1320_ VPWR VGND sg13g2_mux2_1
X_3252_ _1255_ _1257_ _1250_ _1258_ VPWR VGND sg13g2_nand3_1
X_3183_ _1217_ VPWR _0210_ VGND net711 _1166_ sg13g2_o21ai_1
X_2203_ _2022_ _0433_ _0434_ _0435_ VPWR VGND sg13g2_nor3_1
X_2134_ VPWR _1990_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[42\]
+ VGND sg13g2_inv_1
X_2065_ VPWR _1922_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\]
+ VGND sg13g2_inv_1
XFILLER_34_240 VPWR VGND sg13g2_fill_2
XFILLER_34_273 VPWR VGND sg13g2_fill_2
X_2967_ _1090_ VPWR _0120_ VGND net619 _1091_ sg13g2_o21ai_1
X_2898_ _1049_ net78 _1037_ VPWR VGND sg13g2_nand2_1
Xhold620 _0061_ VPWR VGND net939 sg13g2_dlygate4sd3_1
Xhold642 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[3\] VPWR VGND net961 sg13g2_dlygate4sd3_1
Xhold653 u_usb_cdc.endp\[2\] VPWR VGND net972 sg13g2_dlygate4sd3_1
XFILLER_2_829 VPWR VGND sg13g2_decap_8
Xhold631 _0017_ VPWR VGND net950 sg13g2_dlygate4sd3_1
XFILLER_1_339 VPWR VGND sg13g2_decap_8
X_3519_ net972 net766 net587 _0305_ VPWR VGND sg13g2_mux2_1
X_4499_ net701 VGND VPWR _0416_ u_usb_cdc.u_sie.u_phy_tx.data_q\[6\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
Xhold686 u_usb_cdc.u_sie.data_q\[3\] VPWR VGND net1005 sg13g2_dlygate4sd3_1
Xhold675 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] VPWR VGND
+ net994 sg13g2_dlygate4sd3_1
Xhold697 _0260_ VPWR VGND net1016 sg13g2_dlygate4sd3_1
Xhold664 _0373_ VPWR VGND net983 sg13g2_dlygate4sd3_1
XFILLER_40_1006 VPWR VGND sg13g2_decap_8
XFILLER_45_527 VPWR VGND sg13g2_decap_8
XFILLER_27_77 VPWR VGND sg13g2_decap_8
XFILLER_38_590 VPWR VGND sg13g2_fill_2
XFILLER_25_240 VPWR VGND sg13g2_fill_1
XFILLER_40_298 VPWR VGND sg13g2_decap_4
XFILLER_4_15 VPWR VGND sg13g2_decap_4
XFILLER_49_800 VPWR VGND sg13g2_decap_8
XFILLER_0_372 VPWR VGND sg13g2_decap_8
XFILLER_1_884 VPWR VGND sg13g2_decap_8
XFILLER_49_877 VPWR VGND sg13g2_decap_8
XFILLER_36_527 VPWR VGND sg13g2_decap_8
XFILLER_16_284 VPWR VGND sg13g2_fill_1
XFILLER_16_262 VPWR VGND sg13g2_fill_2
XFILLER_20_917 VPWR VGND sg13g2_fill_1
X_3870_ u_usb_cdc.u_sie.u_phy_rx.state_q\[1\] u_usb_cdc.u_sie.u_phy_rx.state_q\[2\]
+ _1744_ _1745_ VPWR VGND sg13g2_nor3_2
X_2821_ VGND VPWR _0994_ _0995_ _0070_ net857 sg13g2_a21oi_1
X_2752_ _0939_ net452 net47 VPWR VGND sg13g2_xnor2_1
XFILLER_9_995 VPWR VGND sg13g2_decap_8
X_2683_ u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\] net57 _0884_ VPWR VGND u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[0\]
+ sg13g2_nand3b_1
X_4422_ net684 VGND VPWR _0350_ u_usb_cdc.sie_out_data\[3\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_2
X_4353_ net676 VGND VPWR net436 u_usb_cdc.u_ctrl_endp.addr_dd\[6\] clknet_leaf_47_clk_regs
+ sg13g2_dfrbpq_1
X_4284_ net650 VGND VPWR net235 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[46\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
X_3304_ VGND VPWR _2008_ net616 _0244_ _1304_ sg13g2_a21oi_1
X_3235_ _1245_ net50 _1156_ VPWR VGND sg13g2_nand2_1
X_3166_ _1208_ VPWR _0202_ VGND _1184_ net609 sg13g2_o21ai_1
X_3097_ _1163_ VPWR _0177_ VGND net828 _1164_ sg13g2_o21ai_1
X_2117_ _1974_ net504 VPWR VGND sg13g2_inv_2
XFILLER_27_549 VPWR VGND sg13g2_decap_8
XFILLER_35_582 VPWR VGND sg13g2_decap_8
XFILLER_23_744 VPWR VGND sg13g2_fill_1
X_3999_ _1833_ net709 _0926_ VPWR VGND sg13g2_nand2_1
XFILLER_13_57 VPWR VGND sg13g2_fill_1
Xhold450 _0286_ VPWR VGND net493 sg13g2_dlygate4sd3_1
Xhold461 u_usb_cdc.u_sie.phy_state_q\[3\] VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold472 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[24\] VPWR VGND
+ net515 sg13g2_dlygate4sd3_1
Xhold494 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[26\] VPWR VGND
+ net537 sg13g2_dlygate4sd3_1
Xhold483 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[6\] VPWR VGND
+ net526 sg13g2_dlygate4sd3_1
XFILLER_49_118 VPWR VGND sg13g2_decap_8
XFILLER_46_869 VPWR VGND sg13g2_decap_8
XFILLER_14_711 VPWR VGND sg13g2_decap_8
XFILLER_14_766 VPWR VGND sg13g2_fill_2
XFILLER_6_965 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_1_692 VPWR VGND sg13g2_decap_8
X_3020_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\] _1019_ net740
+ _1118_ VPWR VGND sg13g2_nand3_1
XFILLER_48_162 VPWR VGND sg13g2_fill_1
XFILLER_49_674 VPWR VGND sg13g2_decap_8
X_3922_ net615 VPWR _1784_ VGND net319 _1780_ sg13g2_o21ai_1
X_3853_ _1733_ VPWR _0364_ VGND _1948_ net595 sg13g2_o21ai_1
X_2804_ _0949_ _0979_ net593 _0980_ VPWR VGND sg13g2_nand3_1
X_3784_ _1682_ VPWR _1683_ VGND net800 _1680_ sg13g2_o21ai_1
X_2735_ _0927_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] _0923_ VPWR VGND sg13g2_nand2_1
X_2666_ _0873_ net844 net596 VPWR VGND sg13g2_nand2_1
X_4405_ net700 VGND VPWR net855 u_usb_cdc.u_sie.crc16_q\[10\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
X_2597_ _0815_ VPWR _0001_ VGND _0720_ _0816_ sg13g2_o21ai_1
X_4336_ net685 VGND VPWR _0264_ u_usb_cdc.u_ctrl_endp.endp_q\[1\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_8_1006 VPWR VGND sg13g2_decap_8
X_4267_ net672 VGND VPWR net273 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[29\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_3218_ _1236_ VPWR _0226_ VGND net720 net603 sg13g2_o21ai_1
X_4198_ net662 VGND VPWR net91 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[44\]
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
X_3149_ _1199_ VPWR _0194_ VGND net720 net607 sg13g2_o21ai_1
XFILLER_11_725 VPWR VGND sg13g2_decap_4
XFILLER_24_89 VPWR VGND sg13g2_fill_2
XFILLER_6_217 VPWR VGND sg13g2_fill_2
XFILLER_40_99 VPWR VGND sg13g2_fill_1
XFILLER_46_1023 VPWR VGND sg13g2_decap_4
Xhold280 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[61\] VPWR
+ VGND net323 sg13g2_dlygate4sd3_1
XFILLER_3_968 VPWR VGND sg13g2_decap_8
Xhold291 _1191_ VPWR VGND net334 sg13g2_dlygate4sd3_1
Xfanout760 net1033 net760 VPWR VGND sg13g2_buf_8
XFILLER_49_75 VPWR VGND sg13g2_decap_8
Xfanout771 u_usb_cdc.bulk_out_nak[0] net771 VPWR VGND sg13g2_buf_8
Xfanout793 net1011 net793 VPWR VGND sg13g2_buf_8
Xfanout782 net783 net782 VPWR VGND sg13g2_buf_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_46_655 VPWR VGND sg13g2_decap_8
XFILLER_14_541 VPWR VGND sg13g2_fill_1
XFILLER_14_552 VPWR VGND sg13g2_decap_4
XFILLER_14_585 VPWR VGND sg13g2_fill_1
XFILLER_41_393 VPWR VGND sg13g2_fill_2
X_2520_ u_usb_cdc.u_ctrl_endp.req_q\[6\] net851 _0747_ VPWR VGND sg13g2_nor2_1
X_2451_ VPWR VGND _0613_ net591 _0610_ net756 _0681_ _0606_ sg13g2_a221oi_1
XFILLER_5_283 VPWR VGND sg13g2_fill_2
X_2382_ u_usb_cdc.u_sie.pid_q\[3\] _0451_ net1053 _0613_ VPWR VGND _0606_ sg13g2_nand4_1
X_4121_ net687 VGND VPWR _0022_ u_usb_cdc.u_sie.phy_state_q\[3\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
X_4052_ _1877_ _1878_ net626 _1880_ VPWR VGND _1879_ sg13g2_nand4_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
X_3003_ _1113_ net135 _1108_ VPWR VGND sg13g2_nand2_1
XFILLER_49_471 VPWR VGND sg13g2_decap_8
X_3905_ _1771_ net714 net391 VPWR VGND sg13g2_nand2_1
X_3836_ _0510_ _0956_ _1722_ VPWR VGND sg13g2_nor2_1
X_3767_ _1667_ _1664_ _1666_ VPWR VGND sg13g2_nand2_1
X_2718_ _0915_ net314 net707 VPWR VGND sg13g2_nand2_1
X_3698_ net777 _0658_ _1601_ VPWR VGND sg13g2_nor2_1
X_2649_ _0860_ u_usb_cdc.u_sie.data_q\[3\] u_usb_cdc.u_sie.data_q\[7\] VPWR VGND sg13g2_xnor2_1
XFILLER_0_916 VPWR VGND sg13g2_decap_8
X_4319_ net651 VGND VPWR net245 net24 clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_25_clk_regs clknet_3_6__leaf_clk_regs clknet_leaf_25_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_28_633 VPWR VGND sg13g2_fill_1
XFILLER_35_44 VPWR VGND sg13g2_fill_1
XFILLER_2_275 VPWR VGND sg13g2_fill_1
Xfanout590 _0618_ net590 VPWR VGND sg13g2_buf_8
XFILLER_47_964 VPWR VGND sg13g2_decap_8
XFILLER_46_474 VPWR VGND sg13g2_decap_4
X_3621_ VGND VPWR net810 _1988_ _1527_ net801 sg13g2_a21oi_1
X_3552_ _1480_ net430 net354 VPWR VGND sg13g2_xnor2_1
X_2503_ _0730_ _0728_ _0729_ _0726_ net623 VPWR VGND sg13g2_a22oi_1
X_3483_ u_usb_cdc.sie_out_data\[6\] _1421_ _1434_ VPWR VGND sg13g2_nor2_1
X_2434_ VGND VPWR _0635_ _0662_ _0664_ _0663_ sg13g2_a21oi_1
X_2365_ _0595_ VPWR _0596_ VGND u_usb_cdc.u_ctrl_endp.state_q\[1\] u_usb_cdc.u_ctrl_endp.state_q\[5\]
+ sg13g2_o21ai_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_4104_ net691 VGND VPWR net412 u_usb_cdc.u_ctrl_endp.req_q\[10\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_2296_ net793 u_usb_cdc.u_ctrl_endp.max_length_q\[0\] _0528_ VPWR VGND sg13g2_xor2_1
X_4035_ _1865_ net356 net642 VPWR VGND sg13g2_nand2_1
XFILLER_36_1000 VPWR VGND sg13g2_decap_8
X_3819_ _1708_ _0973_ _1701_ VPWR VGND sg13g2_nand2_1
XFILLER_21_46 VPWR VGND sg13g2_fill_2
XFILLER_0_713 VPWR VGND sg13g2_decap_8
XFILLER_48_717 VPWR VGND sg13g2_decap_8
XFILLER_29_931 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_fill_2
XFILLER_44_956 VPWR VGND sg13g2_decap_8
XFILLER_24_691 VPWR VGND sg13g2_fill_1
XFILLER_7_378 VPWR VGND sg13g2_fill_1
XFILLER_7_389 VPWR VGND sg13g2_decap_4
X_2150_ VPWR _2006_ net174 VGND sg13g2_inv_1
X_2081_ VPWR _1938_ net794 VGND sg13g2_inv_1
XFILLER_47_761 VPWR VGND sg13g2_decap_8
XFILLER_35_934 VPWR VGND sg13g2_fill_2
X_2983_ _1102_ VPWR _0125_ VGND _1048_ net610 sg13g2_o21ai_1
X_3604_ _1510_ _0541_ _0655_ VPWR VGND sg13g2_nand2b_1
X_3535_ u_usb_cdc.u_ctrl_endp.addr_dd\[2\] u_usb_cdc.u_ctrl_endp.addr_dd\[5\] u_usb_cdc.u_ctrl_endp.addr_dd\[4\]
+ u_usb_cdc.u_ctrl_endp.addr_dd\[6\] _1467_ VPWR VGND sg13g2_nor4_1
X_3466_ VGND VPWR net576 _1422_ _0288_ _1420_ sg13g2_a21oi_1
X_2417_ net782 net784 _0647_ VPWR VGND sg13g2_nor2b_2
X_3397_ _1381_ _1379_ _1380_ VPWR VGND sg13g2_nand2_1
X_2348_ net836 net837 _0577_ _0579_ _0580_ VPWR VGND sg13g2_nor4_1
X_2279_ VPWR _0511_ _0510_ VGND sg13g2_inv_1
X_4018_ _1850_ _1967_ u_usb_cdc.u_sie.phy_state_q\[10\] u_usb_cdc.u_sie.data_q\[3\]
+ net842 VPWR VGND sg13g2_a22oi_1
XFILLER_26_967 VPWR VGND sg13g2_decap_8
XFILLER_37_271 VPWR VGND sg13g2_decap_4
XFILLER_13_639 VPWR VGND sg13g2_fill_1
XFILLER_32_23 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_40_clk_regs clknet_3_5__leaf_clk_regs clknet_leaf_40_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_0_554 VPWR VGND sg13g2_decap_8
XFILLER_0_598 VPWR VGND sg13g2_fill_1
XFILLER_17_901 VPWR VGND sg13g2_decap_8
XFILLER_44_720 VPWR VGND sg13g2_decap_8
XFILLER_32_904 VPWR VGND sg13g2_decap_8
XFILLER_44_753 VPWR VGND sg13g2_decap_8
XFILLER_8_610 VPWR VGND sg13g2_decap_8
XFILLER_12_661 VPWR VGND sg13g2_fill_1
XFILLER_40_992 VPWR VGND sg13g2_decap_8
XFILLER_8_665 VPWR VGND sg13g2_fill_2
XFILLER_8_698 VPWR VGND sg13g2_fill_2
Xhold109 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[64\] VPWR
+ VGND net152 sg13g2_dlygate4sd3_1
Xheichips25_usb_cdc_41 VPWR VGND uio_oe[5] sg13g2_tiehi
X_3320_ _1318_ VPWR _1319_ VGND net818 net125 sg13g2_o21ai_1
X_3251_ _1257_ net813 _1256_ VPWR VGND sg13g2_xnor2_1
X_3182_ _1217_ net127 _1213_ VPWR VGND sg13g2_nand2_1
X_2202_ _0434_ _1921_ net368 VPWR VGND sg13g2_nand2_1
XFILLER_39_503 VPWR VGND sg13g2_fill_2
X_2133_ VPWR _1989_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[41\]
+ VGND sg13g2_inv_1
X_2064_ VPWR _1921_ net835 VGND sg13g2_inv_1
XFILLER_31_981 VPWR VGND sg13g2_decap_8
X_2966_ _1091_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2897_ _1047_ VPWR _0093_ VGND net618 _1048_ sg13g2_o21ai_1
Xhold621 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[2\] VPWR VGND
+ net940 sg13g2_dlygate4sd3_1
Xhold610 u_usb_cdc.u_sie.u_phy_rx.state_q\[3\] VPWR VGND net929 sg13g2_dlygate4sd3_1
Xhold643 _1740_ VPWR VGND net962 sg13g2_dlygate4sd3_1
Xhold654 u_usb_cdc.u_sie.crc16_q\[4\] VPWR VGND net973 sg13g2_dlygate4sd3_1
Xhold632 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[3\] VPWR VGND
+ net951 sg13g2_dlygate4sd3_1
X_3518_ net995 net767 net587 _0304_ VPWR VGND sg13g2_mux2_1
Xhold676 u_usb_cdc.endp\[1\] VPWR VGND net995 sg13g2_dlygate4sd3_1
XFILLER_1_318 VPWR VGND sg13g2_decap_8
X_4498_ net701 VGND VPWR net357 u_usb_cdc.u_sie.u_phy_tx.data_q\[5\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
Xhold687 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ VPWR VGND net1006 sg13g2_dlygate4sd3_1
Xhold665 u_usb_cdc.u_sie.data_q\[7\] VPWR VGND net984 sg13g2_dlygate4sd3_1
X_3449_ _0283_ _1410_ net179 VPWR VGND sg13g2_nand2b_1
Xhold698 u_usb_cdc.u_sie.phy_state_q\[8\] VPWR VGND net1017 sg13g2_dlygate4sd3_1
XFILLER_17_208 VPWR VGND sg13g2_fill_2
XFILLER_27_56 VPWR VGND sg13g2_decap_8
XFILLER_26_764 VPWR VGND sg13g2_fill_2
XFILLER_14_948 VPWR VGND sg13g2_fill_1
XFILLER_40_233 VPWR VGND sg13g2_fill_2
XFILLER_40_222 VPWR VGND sg13g2_fill_2
XFILLER_49_1010 VPWR VGND sg13g2_decap_8
XFILLER_0_351 VPWR VGND sg13g2_decap_8
XFILLER_49_856 VPWR VGND sg13g2_decap_8
XFILLER_48_366 VPWR VGND sg13g2_fill_1
XFILLER_36_517 VPWR VGND sg13g2_fill_1
XFILLER_31_222 VPWR VGND sg13g2_fill_1
XFILLER_32_745 VPWR VGND sg13g2_fill_2
X_2820_ net742 _0961_ _0995_ VPWR VGND sg13g2_and2_1
X_2751_ _0938_ net532 net48 VPWR VGND sg13g2_xnor2_1
X_2682_ _2036_ _0882_ _0883_ VPWR VGND sg13g2_nor2_1
XFILLER_9_974 VPWR VGND sg13g2_decap_8
X_4421_ net684 VGND VPWR _0349_ u_usb_cdc.sie_out_data\[2\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_2
X_4352_ net676 VGND VPWR net474 u_usb_cdc.u_ctrl_endp.addr_dd\[5\] clknet_leaf_47_clk_regs
+ sg13g2_dfrbpq_1
X_4283_ net655 VGND VPWR net163 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[45\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_3303_ VPWR VGND _1983_ net616 _1303_ net129 _1304_ net629 sg13g2_a221oi_1
X_3234_ _1244_ VPWR _0234_ VGND _1155_ _1184_ sg13g2_o21ai_1
X_3165_ _1208_ net125 net609 VPWR VGND sg13g2_nand2_1
X_3096_ net832 _1159_ net761 _1164_ VPWR VGND sg13g2_nand3_1
X_2116_ VPWR _1973_ net301 VGND sg13g2_inv_1
XFILLER_35_550 VPWR VGND sg13g2_fill_2
XFILLER_23_723 VPWR VGND sg13g2_decap_8
XFILLER_10_406 VPWR VGND sg13g2_decap_4
X_3998_ _2027_ _0925_ _1832_ VPWR VGND sg13g2_nor2_1
X_2949_ _1079_ net636 VPWR VGND net620 sg13g2_nand2b_2
Xhold440 u_usb_cdc.u_ctrl_endp.req_q\[6\] VPWR VGND net483 sg13g2_dlygate4sd3_1
Xhold462 _0028_ VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold451 u_usb_cdc.u_sie.u_phy_tx.data_q\[6\] VPWR VGND net494 sg13g2_dlygate4sd3_1
Xhold495 _0109_ VPWR VGND net538 sg13g2_dlygate4sd3_1
Xhold473 _0107_ VPWR VGND net516 sg13g2_dlygate4sd3_1
Xhold484 _0089_ VPWR VGND net527 sg13g2_dlygate4sd3_1
XFILLER_38_11 VPWR VGND sg13g2_decap_4
XFILLER_38_44 VPWR VGND sg13g2_decap_4
XFILLER_46_848 VPWR VGND sg13g2_decap_8
XFILLER_45_347 VPWR VGND sg13g2_fill_1
XFILLER_26_583 VPWR VGND sg13g2_fill_2
XFILLER_14_756 VPWR VGND sg13g2_fill_1
XFILLER_41_586 VPWR VGND sg13g2_fill_1
XFILLER_10_973 VPWR VGND sg13g2_decap_8
XFILLER_5_487 VPWR VGND sg13g2_decap_8
XFILLER_1_671 VPWR VGND sg13g2_decap_8
XFILLER_23_1013 VPWR VGND sg13g2_decap_8
XFILLER_49_653 VPWR VGND sg13g2_decap_8
XFILLER_37_859 VPWR VGND sg13g2_fill_2
X_3921_ net319 _1780_ _1783_ VPWR VGND sg13g2_and2_1
X_3852_ _0899_ _1729_ net329 _1733_ VPWR VGND sg13g2_nand3_1
X_2803_ VGND VPWR net844 _0978_ _0979_ _0976_ sg13g2_a21oi_1
XFILLER_30_1017 VPWR VGND sg13g2_decap_8
X_3783_ VGND VPWR net800 _1681_ _1682_ _1923_ sg13g2_a21oi_1
X_2734_ VPWR VGND _1979_ _0925_ _0923_ net625 _0036_ _2028_ sg13g2_a221oi_1
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
X_2665_ _0024_ _0872_ _1973_ _0599_ net601 VPWR VGND sg13g2_a22oi_1
X_2596_ _0707_ _0727_ _0729_ _0816_ VPWR VGND sg13g2_or3_1
X_4404_ net696 VGND VPWR net889 u_usb_cdc.u_sie.crc16_q\[9\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
X_4335_ net683 VGND VPWR _0263_ u_usb_cdc.u_ctrl_endp.endp_q\[0\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
X_4266_ net654 VGND VPWR net281 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[28\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_3217_ _1236_ net211 net603 VPWR VGND sg13g2_nand2_1
X_4197_ net662 VGND VPWR net60 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[43\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
X_3148_ _1199_ net195 net607 VPWR VGND sg13g2_nand2_1
X_3079_ _1150_ net202 net635 VPWR VGND sg13g2_nand2_1
XFILLER_3_914 VPWR VGND sg13g2_decap_4
XFILLER_3_947 VPWR VGND sg13g2_decap_8
XFILLER_46_1002 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_fill_1
Xhold270 _0361_ VPWR VGND net313 sg13g2_dlygate4sd3_1
Xhold281 _0228_ VPWR VGND net324 sg13g2_dlygate4sd3_1
Xhold292 _0190_ VPWR VGND net335 sg13g2_dlygate4sd3_1
XFILLER_49_54 VPWR VGND sg13g2_decap_8
Xfanout750 net751 net750 VPWR VGND sg13g2_buf_8
Xfanout794 net946 net794 VPWR VGND sg13g2_buf_8
Xfanout761 net1045 net761 VPWR VGND sg13g2_buf_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
Xfanout772 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] net772 VPWR VGND sg13g2_buf_8
Xfanout783 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[3\] net783 VPWR VGND sg13g2_buf_2
X_2450_ VPWR VGND _0644_ net590 net588 net756 _0680_ _0606_ sg13g2_a221oi_1
X_2381_ _0612_ net755 _0606_ VPWR VGND sg13g2_nand2_2
XFILLER_39_4 VPWR VGND sg13g2_decap_8
X_4120_ net687 VGND VPWR net525 u_usb_cdc.u_sie.phy_state_q\[2\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
X_4051_ _1879_ _1962_ net837 u_usb_cdc.u_sie.data_q\[7\] net843 VPWR VGND sg13g2_a22oi_1
XFILLER_49_450 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
X_3002_ _1112_ VPWR _0134_ VGND _1068_ net610 sg13g2_o21ai_1
X_3904_ _1768_ VPWR _0378_ VGND _1769_ _1770_ sg13g2_o21ai_1
X_3835_ net756 VPWR _1721_ VGND _1719_ _1720_ sg13g2_o21ai_1
XFILLER_20_578 VPWR VGND sg13g2_fill_2
X_3766_ VGND VPWR net800 _1665_ _1666_ _1923_ sg13g2_a21oi_1
X_2717_ _0031_ _0912_ _0914_ VPWR VGND sg13g2_nand2_1
X_3697_ _1520_ _1543_ _0653_ _1600_ VPWR VGND sg13g2_nand3_1
X_2648_ _0859_ net766 u_usb_cdc.u_sie.data_q\[5\] VPWR VGND sg13g2_xnor2_1
X_2579_ _0803_ net719 _0641_ VPWR VGND sg13g2_nand2_1
X_4318_ net648 VGND VPWR net52 net23 clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
X_4249_ net649 VGND VPWR net279 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[11\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
XFILLER_19_68 VPWR VGND sg13g2_fill_2
XFILLER_28_667 VPWR VGND sg13g2_fill_2
XFILLER_43_637 VPWR VGND sg13g2_fill_2
XFILLER_7_505 VPWR VGND sg13g2_fill_1
Xfanout580 _1493_ net580 VPWR VGND sg13g2_buf_8
Xfanout591 _0618_ net591 VPWR VGND sg13g2_buf_2
XFILLER_47_943 VPWR VGND sg13g2_decap_8
XFILLER_18_133 VPWR VGND sg13g2_decap_4
XFILLER_19_645 VPWR VGND sg13g2_fill_2
XFILLER_34_637 VPWR VGND sg13g2_fill_1
X_3620_ net810 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[0\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[8\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[16\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[24\]
+ net801 _1526_ VPWR VGND sg13g2_mux4_1
X_3551_ _1479_ net430 _1476_ VPWR VGND sg13g2_nand2_1
X_2502_ _1937_ net794 u_usb_cdc.u_ctrl_endp.rec_q\[0\] _0729_ VPWR VGND u_usb_cdc.configured_o
+ sg13g2_nand4_1
X_3482_ net564 net577 _1433_ VPWR VGND sg13g2_nor2_1
X_2433_ net590 _0621_ net624 _0661_ _0663_ VPWR VGND sg13g2_nor4_1
X_2364_ _0595_ u_usb_cdc.sie_in_req net640 VPWR VGND sg13g2_nand2_2
X_4103_ net691 VGND VPWR _0010_ u_usb_cdc.u_ctrl_endp.req_q\[9\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_2295_ u_usb_cdc.u_ctrl_endp.max_length_q\[4\] net778 _0527_ VPWR VGND sg13g2_xor2_1
X_4034_ _1858_ VPWR _0414_ VGND _1863_ _1864_ sg13g2_o21ai_1
XFILLER_21_821 VPWR VGND sg13g2_decap_8
XFILLER_32_180 VPWR VGND sg13g2_fill_1
X_3818_ _1707_ net911 _1703_ _0355_ VPWR VGND sg13g2_mux2_1
X_3749_ _1643_ VPWR _1650_ VGND _1646_ _1649_ sg13g2_o21ai_1
XFILLER_0_769 VPWR VGND sg13g2_decap_8
XFILLER_46_33 VPWR VGND sg13g2_decap_8
XFILLER_29_987 VPWR VGND sg13g2_decap_8
XFILLER_46_66 VPWR VGND sg13g2_fill_2
XFILLER_44_935 VPWR VGND sg13g2_decap_8
XFILLER_11_342 VPWR VGND sg13g2_decap_8
XFILLER_8_869 VPWR VGND sg13g2_decap_8
X_2080_ VPWR _1937_ u_usb_cdc.u_ctrl_endp.rec_q\[1\] VGND sg13g2_inv_1
XFILLER_47_740 VPWR VGND sg13g2_decap_8
XFILLER_46_250 VPWR VGND sg13g2_fill_2
XFILLER_19_486 VPWR VGND sg13g2_fill_1
X_2982_ _1102_ net74 _1096_ VPWR VGND sg13g2_nand2_1
XFILLER_22_618 VPWR VGND sg13g2_decap_8
XFILLER_21_128 VPWR VGND sg13g2_fill_1
X_3603_ VGND VPWR _1506_ _1508_ _1509_ _0537_ sg13g2_a21oi_1
X_3534_ _1466_ _0619_ _1465_ u_usb_cdc.bus_reset net742 VPWR VGND sg13g2_a22oi_1
X_3465_ net763 _1421_ _1422_ VPWR VGND sg13g2_nor2_1
X_2416_ VPWR _0646_ _0645_ VGND sg13g2_inv_1
X_3396_ net802 net809 net797 _1380_ VPWR VGND sg13g2_a21o_1
X_2347_ net710 _0578_ _0579_ VPWR VGND sg13g2_nor2_1
X_2278_ _0498_ _0509_ _0497_ _0510_ VPWR VGND sg13g2_nand3_1
X_4017_ _1849_ _1956_ net845 u_usb_cdc.u_sie.pid_q\[3\] net836 VPWR VGND sg13g2_a22oi_1
XFILLER_41_949 VPWR VGND sg13g2_decap_8
XFILLER_12_117 VPWR VGND sg13g2_fill_2
XFILLER_32_35 VPWR VGND sg13g2_decap_4
XFILLER_5_817 VPWR VGND sg13g2_fill_1
XFILLER_5_839 VPWR VGND sg13g2_fill_2
XFILLER_10_1004 VPWR VGND sg13g2_decap_8
XFILLER_0_533 VPWR VGND sg13g2_decap_8
XFILLER_48_559 VPWR VGND sg13g2_fill_1
XFILLER_17_946 VPWR VGND sg13g2_fill_2
XFILLER_25_990 VPWR VGND sg13g2_decap_8
XFILLER_40_971 VPWR VGND sg13g2_decap_8
XFILLER_12_673 VPWR VGND sg13g2_fill_1
Xheichips25_usb_cdc_42 VPWR VGND uio_oe[6] sg13g2_tiehi
X_3250_ _1256_ net827 _1193_ VPWR VGND sg13g2_xnor2_1
X_3181_ _1216_ VPWR _0209_ VGND net712 _1164_ sg13g2_o21ai_1
X_2201_ _0433_ net626 net709 VPWR VGND sg13g2_nand2_1
X_2132_ VPWR _1988_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[40\]
+ VGND sg13g2_inv_1
X_2063_ VPWR _1920_ net836 VGND sg13g2_inv_1
XFILLER_34_275 VPWR VGND sg13g2_fill_1
XFILLER_31_960 VPWR VGND sg13g2_decap_8
X_2965_ _1090_ net113 _1079_ VPWR VGND sg13g2_nand2_1
X_2896_ _1048_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net645 VPWR VGND sg13g2_nand2_1
Xhold600 _0391_ VPWR VGND net919 sg13g2_dlygate4sd3_1
Xhold611 _0035_ VPWR VGND net930 sg13g2_dlygate4sd3_1
Xhold644 _1741_ VPWR VGND net963 sg13g2_dlygate4sd3_1
X_3517_ VGND VPWR net719 net586 _0303_ _1458_ sg13g2_a21oi_1
Xhold633 _0254_ VPWR VGND net952 sg13g2_dlygate4sd3_1
Xhold622 _0253_ VPWR VGND net941 sg13g2_dlygate4sd3_1
Xhold688 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] VPWR VGND net1007 sg13g2_dlygate4sd3_1
Xhold666 net19 VPWR VGND net985 sg13g2_dlygate4sd3_1
X_4497_ net701 VGND VPWR net293 u_usb_cdc.u_sie.u_phy_tx.data_q\[4\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
Xhold655 u_usb_cdc.u_ctrl_endp.req_q\[8\] VPWR VGND net974 sg13g2_dlygate4sd3_1
Xhold677 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ VPWR VGND net996 sg13g2_dlygate4sd3_1
X_3448_ net623 net489 _1410_ _0282_ VPWR VGND sg13g2_mux2_1
Xhold699 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ VPWR VGND net1018 sg13g2_dlygate4sd3_1
X_3379_ net629 _1365_ _1366_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_35 VPWR VGND sg13g2_decap_8
XFILLER_38_592 VPWR VGND sg13g2_fill_1
XFILLER_43_67 VPWR VGND sg13g2_fill_2
XFILLER_1_820 VPWR VGND sg13g2_fill_1
XFILLER_0_330 VPWR VGND sg13g2_decap_8
XFILLER_49_835 VPWR VGND sg13g2_decap_8
XFILLER_48_334 VPWR VGND sg13g2_fill_1
XFILLER_1_1024 VPWR VGND sg13g2_decap_4
XFILLER_17_743 VPWR VGND sg13g2_fill_2
XFILLER_32_757 VPWR VGND sg13g2_fill_1
XFILLER_9_953 VPWR VGND sg13g2_fill_1
X_2750_ _0042_ _0936_ _0937_ VPWR VGND sg13g2_nand2_1
X_2681_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\] u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[0\]
+ _0882_ VPWR VGND sg13g2_nor2_1
X_4420_ net684 VGND VPWR _0348_ u_usb_cdc.sie_out_data\[1\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_8_496 VPWR VGND sg13g2_decap_8
X_4351_ net676 VGND VPWR _0279_ u_usb_cdc.u_ctrl_endp.addr_dd\[4\] clknet_leaf_51_clk_regs
+ sg13g2_dfrbpq_1
X_3302_ _1302_ VPWR _1303_ VGND _1286_ _1300_ sg13g2_o21ai_1
X_4282_ net655 VGND VPWR net231 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[44\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_3233_ _1244_ net191 _1156_ VPWR VGND sg13g2_nand2_1
X_3164_ _1207_ VPWR _0201_ VGND _1182_ net608 sg13g2_o21ai_1
XFILLER_12_0 VPWR VGND sg13g2_fill_2
X_3095_ _1163_ net66 _1151_ VPWR VGND sg13g2_nand2_1
X_2115_ _1972_ net921 VPWR VGND sg13g2_inv_2
X_3997_ _0410_ _1829_ _1831_ net643 _1993_ VPWR VGND sg13g2_a22oi_1
X_2948_ _1034_ _1018_ _1078_ VPWR VGND sg13g2_nor2b_2
X_2879_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net443 _1036_ _0087_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_19_clk_regs clknet_3_3__leaf_clk_regs clknet_leaf_19_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_2_639 VPWR VGND sg13g2_decap_8
Xhold441 _0007_ VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold430 u_usb_cdc.u_ctrl_endp.addr_dd\[5\] VPWR VGND net473 sg13g2_dlygate4sd3_1
XFILLER_8_8 VPWR VGND sg13g2_fill_2
Xhold452 _1876_ VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold463 u_usb_cdc.u_sie.rx_data\[6\] VPWR VGND net506 sg13g2_dlygate4sd3_1
Xhold496 u_usb_cdc.u_sie.crc16_q\[5\] VPWR VGND net539 sg13g2_dlygate4sd3_1
Xhold474 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[57\] VPWR VGND
+ net517 sg13g2_dlygate4sd3_1
Xhold485 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[27\] VPWR VGND
+ net528 sg13g2_dlygate4sd3_1
XFILLER_46_816 VPWR VGND sg13g2_decap_4
XFILLER_46_827 VPWR VGND sg13g2_decap_8
XFILLER_14_779 VPWR VGND sg13g2_fill_1
XFILLER_5_466 VPWR VGND sg13g2_decap_8
XFILLER_1_650 VPWR VGND sg13g2_decap_8
XFILLER_0_171 VPWR VGND sg13g2_decap_4
XFILLER_49_632 VPWR VGND sg13g2_decap_8
XFILLER_37_838 VPWR VGND sg13g2_fill_1
XFILLER_17_540 VPWR VGND sg13g2_fill_2
XFILLER_17_573 VPWR VGND sg13g2_decap_8
X_3920_ _1782_ net713 net319 VPWR VGND sg13g2_nand2_1
X_3851_ _1732_ VPWR _0363_ VGND _1949_ net595 sg13g2_o21ai_1
X_2802_ _0978_ _0974_ _0977_ VPWR VGND sg13g2_nand2_1
XFILLER_32_587 VPWR VGND sg13g2_fill_2
XFILLER_20_738 VPWR VGND sg13g2_decap_4
X_3782_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[55\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[63\]
+ net808 _1681_ VPWR VGND sg13g2_mux2_1
XFILLER_9_750 VPWR VGND sg13g2_fill_1
X_2733_ VGND VPWR _0926_ u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\]
+ sg13g2_or2_1
X_2664_ net601 VPWR _0872_ VGND net838 _0871_ sg13g2_o21ai_1
X_2595_ net522 VPWR _0815_ VGND _0812_ _0814_ sg13g2_o21ai_1
X_4403_ net696 VGND VPWR net916 u_usb_cdc.u_sie.crc16_q\[8\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
X_4334_ net682 VGND VPWR net981 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\]
+ clknet_leaf_20_clk_regs sg13g2_dfrbpq_2
X_4265_ net656 VGND VPWR _0194_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[27\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_3216_ _1235_ VPWR _0225_ VGND _1913_ net603 sg13g2_o21ai_1
X_4196_ net660 VGND VPWR net75 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[42\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
X_3147_ VGND VPWR _1995_ net605 _0193_ _1198_ sg13g2_a21oi_1
X_3078_ _1149_ VPWR _0173_ VGND _1917_ net635 sg13g2_o21ai_1
XFILLER_23_532 VPWR VGND sg13g2_fill_1
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_23_576 VPWR VGND sg13g2_decap_4
Xhold271 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[4\] VPWR VGND net314 sg13g2_dlygate4sd3_1
Xhold260 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[60\] VPWR
+ VGND net303 sg13g2_dlygate4sd3_1
Xhold282 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[18\] VPWR
+ VGND net325 sg13g2_dlygate4sd3_1
XFILLER_49_33 VPWR VGND sg13g2_decap_8
Xhold293 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[2\] VPWR VGND net336 sg13g2_dlygate4sd3_1
Xfanout751 net934 net751 VPWR VGND sg13g2_buf_8
Xfanout740 net741 net740 VPWR VGND sg13g2_buf_2
Xfanout762 u_usb_cdc.sie_out_data\[1\] net762 VPWR VGND sg13g2_buf_8
XFILLER_49_99 VPWR VGND sg13g2_fill_1
Xfanout784 net786 net784 VPWR VGND sg13g2_buf_2
Xfanout773 net775 net773 VPWR VGND sg13g2_buf_8
Xfanout795 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\] net795
+ VPWR VGND sg13g2_buf_8
XFILLER_45_145 VPWR VGND sg13g2_fill_1
XFILLER_42_896 VPWR VGND sg13g2_decap_8
XFILLER_6_775 VPWR VGND sg13g2_decap_4
XFILLER_6_797 VPWR VGND sg13g2_decap_4
X_2380_ _0611_ _0609_ VPWR VGND _0598_ sg13g2_nand2b_2
X_4050_ _1878_ _1961_ net845 _1935_ u_usb_cdc.u_sie.phy_state_q\[11\] VPWR VGND sg13g2_a22oi_1
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
X_3001_ _1112_ net86 _1108_ VPWR VGND sg13g2_nand2_1
X_3903_ net615 VPWR _1770_ VGND net457 _1765_ sg13g2_o21ai_1
X_3834_ net840 _0436_ _1474_ _1720_ VPWR VGND sg13g2_nor3_1
X_3765_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[54\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[62\]
+ net808 _1665_ VPWR VGND sg13g2_mux2_1
X_2716_ VGND VPWR net961 net707 _0914_ _0913_ sg13g2_a21oi_1
X_3696_ _1586_ VPWR _1599_ VGND net795 _1598_ sg13g2_o21ai_1
X_2647_ _0858_ net767 u_usb_cdc.u_sie.data_q\[4\] VPWR VGND sg13g2_xnor2_1
X_2578_ _0801_ VPWR _0007_ VGND _0720_ _0802_ sg13g2_o21ai_1
X_4317_ net648 VGND VPWR net447 net22 clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
X_4248_ net654 VGND VPWR net67 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[10\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
XFILLER_28_613 VPWR VGND sg13g2_decap_8
X_4179_ net666 VGND VPWR net512 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[25\]
+ clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
XFILLER_24_896 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_34_clk_regs clknet_3_6__leaf_clk_regs clknet_leaf_34_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_13_1024 VPWR VGND sg13g2_decap_4
XFILLER_47_922 VPWR VGND sg13g2_decap_8
Xfanout592 net594 net592 VPWR VGND sg13g2_buf_8
Xfanout581 _1401_ net581 VPWR VGND sg13g2_buf_8
XFILLER_18_112 VPWR VGND sg13g2_fill_1
XFILLER_46_421 VPWR VGND sg13g2_fill_2
XFILLER_47_999 VPWR VGND sg13g2_decap_8
XFILLER_18_156 VPWR VGND sg13g2_fill_1
XFILLER_33_126 VPWR VGND sg13g2_fill_2
XFILLER_15_841 VPWR VGND sg13g2_fill_1
XFILLER_33_137 VPWR VGND sg13g2_fill_2
XFILLER_42_671 VPWR VGND sg13g2_decap_8
XFILLER_42_682 VPWR VGND sg13g2_fill_1
X_3550_ _1478_ VPWR _0316_ VGND net354 _1477_ sg13g2_o21ai_1
X_2501_ _0707_ _0727_ _0728_ VPWR VGND sg13g2_nor2_1
X_3481_ VGND VPWR net577 _1432_ _0293_ _1431_ sg13g2_a21oi_1
X_2432_ net590 _0621_ net624 _0662_ VPWR VGND sg13g2_nor3_2
X_2363_ VGND VPWR _0592_ _0593_ _0594_ _0516_ sg13g2_a21oi_1
X_4102_ net693 VGND VPWR net975 u_usb_cdc.u_ctrl_endp.req_q\[8\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_2_61 VPWR VGND sg13g2_fill_1
X_4033_ net625 VPWR _1864_ VGND u_usb_cdc.u_sie.u_phy_tx.data_q\[5\] _2026_ sg13g2_o21ai_1
X_2294_ net772 u_usb_cdc.u_ctrl_endp.max_length_q\[6\] _0526_ VPWR VGND sg13g2_xor2_1
XFILLER_38_988 VPWR VGND sg13g2_decap_8
X_3817_ _1707_ _1705_ _1706_ VPWR VGND sg13g2_nand2_1
X_3748_ net796 VPWR _1649_ VGND _1647_ _1648_ sg13g2_o21ai_1
X_3679_ VPWR VGND net637 net627 _1582_ _1499_ _1583_ _1573_ sg13g2_a221oi_1
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_43_1017 VPWR VGND sg13g2_decap_8
XFILLER_0_748 VPWR VGND sg13g2_decap_8
XFILLER_29_966 VPWR VGND sg13g2_decap_8
XFILLER_46_23 VPWR VGND sg13g2_fill_1
XFILLER_47_229 VPWR VGND sg13g2_fill_1
XFILLER_44_914 VPWR VGND sg13g2_decap_8
XFILLER_23_170 VPWR VGND sg13g2_fill_2
XFILLER_12_899 VPWR VGND sg13g2_decap_8
XFILLER_38_229 VPWR VGND sg13g2_fill_2
XFILLER_47_796 VPWR VGND sg13g2_decap_8
XFILLER_15_682 VPWR VGND sg13g2_fill_2
X_2981_ _1101_ VPWR _0124_ VGND _1046_ net610 sg13g2_o21ai_1
XFILLER_30_652 VPWR VGND sg13g2_fill_2
X_3602_ _1508_ _1507_ net782 VPWR VGND sg13g2_nand2b_1
X_3533_ VGND VPWR _1940_ _1396_ _1465_ _0588_ sg13g2_a21oi_1
X_3464_ _0661_ VPWR _1421_ VGND net719 _0751_ sg13g2_o21ai_1
XFILLER_42_0 VPWR VGND sg13g2_decap_4
X_2415_ _0645_ net787 _0634_ VPWR VGND sg13g2_nand2_2
X_3395_ net802 net797 net809 _1379_ VPWR VGND sg13g2_nand3_1
X_2346_ VGND VPWR _0578_ _0510_ _0506_ sg13g2_or2_1
X_2277_ _0488_ _0494_ _0507_ _0508_ _0509_ VPWR VGND sg13g2_nor4_1
X_4016_ net642 net439 _1848_ _0412_ VPWR VGND sg13g2_a21o_1
XFILLER_26_903 VPWR VGND sg13g2_decap_8
XFILLER_41_928 VPWR VGND sg13g2_decap_8
XFILLER_34_980 VPWR VGND sg13g2_decap_8
XFILLER_32_25 VPWR VGND sg13g2_fill_1
XFILLER_20_151 VPWR VGND sg13g2_decap_8
XFILLER_20_162 VPWR VGND sg13g2_fill_1
XFILLER_4_317 VPWR VGND sg13g2_fill_2
XFILLER_0_512 VPWR VGND sg13g2_decap_8
XFILLER_0_589 VPWR VGND sg13g2_decap_8
XFILLER_44_700 VPWR VGND sg13g2_decap_8
XFILLER_28_284 VPWR VGND sg13g2_fill_1
XFILLER_43_243 VPWR VGND sg13g2_decap_4
XFILLER_44_788 VPWR VGND sg13g2_decap_8
XFILLER_40_950 VPWR VGND sg13g2_decap_8
Xheichips25_usb_cdc_32 VPWR VGND uio_oe[0] sg13g2_tielo
Xheichips25_usb_cdc_43 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_3_372 VPWR VGND sg13g2_decap_8
XFILLER_3_350 VPWR VGND sg13g2_fill_2
X_2200_ _2048_ _2049_ _0430_ _0432_ _0064_ VPWR VGND sg13g2_and4_1
XFILLER_26_1023 VPWR VGND sg13g2_decap_4
X_3180_ _1216_ net175 _1213_ VPWR VGND sg13g2_nand2_1
X_2131_ VPWR _1987_ net486 VGND sg13g2_inv_1
X_2062_ _1919_ net843 VPWR VGND sg13g2_inv_2
X_2964_ _1088_ VPWR _0119_ VGND net619 _1089_ sg13g2_o21ai_1
XFILLER_33_1005 VPWR VGND sg13g2_decap_8
X_2895_ _1047_ net76 _1037_ VPWR VGND sg13g2_nand2_1
Xhold601 u_usb_cdc.u_sie.crc16_q\[11\] VPWR VGND net920 sg13g2_dlygate4sd3_1
Xhold612 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[0\] VPWR VGND
+ net931 sg13g2_dlygate4sd3_1
Xhold645 _0368_ VPWR VGND net964 sg13g2_dlygate4sd3_1
Xhold634 u_usb_cdc.u_ctrl_endp.rec_q\[1\] VPWR VGND net953 sg13g2_dlygate4sd3_1
X_3516_ net993 net586 _1458_ VPWR VGND sg13g2_nor2_1
Xhold623 u_usb_cdc.u_ctrl_endp.req_q\[3\] VPWR VGND net942 sg13g2_dlygate4sd3_1
Xhold667 u_usb_cdc.u_sie.phy_state_q\[11\] VPWR VGND net986 sg13g2_dlygate4sd3_1
X_4496_ net701 VGND VPWR net384 u_usb_cdc.u_sie.u_phy_tx.data_q\[3\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
Xhold656 _0009_ VPWR VGND net975 sg13g2_dlygate4sd3_1
Xhold678 u_usb_cdc.u_sie.data_q\[4\] VPWR VGND net997 sg13g2_dlygate4sd3_1
Xhold689 _0030_ VPWR VGND net1008 sg13g2_dlygate4sd3_1
X_3447_ _1388_ VPWR _1410_ VGND _1398_ _1409_ sg13g2_o21ai_1
X_3378_ net814 net813 net820 _1365_ VPWR VGND sg13g2_nand3_1
X_2329_ _0558_ _0560_ u_usb_cdc.endp\[0\] _0561_ VPWR VGND sg13g2_nand3_1
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_25_221 VPWR VGND sg13g2_fill_2
XFILLER_40_235 VPWR VGND sg13g2_fill_1
XFILLER_41_758 VPWR VGND sg13g2_decap_8
XFILLER_41_769 VPWR VGND sg13g2_fill_1
XFILLER_49_814 VPWR VGND sg13g2_decap_8
XFILLER_0_386 VPWR VGND sg13g2_decap_8
XFILLER_1_898 VPWR VGND sg13g2_decap_8
XFILLER_1_1003 VPWR VGND sg13g2_decap_8
XFILLER_44_530 VPWR VGND sg13g2_decap_8
XFILLER_32_736 VPWR VGND sg13g2_decap_4
XFILLER_32_747 VPWR VGND sg13g2_fill_1
X_2680_ _0881_ net1007 _2042_ VPWR VGND sg13g2_nand2_1
X_4350_ net683 VGND VPWR _0278_ u_usb_cdc.u_ctrl_endp.addr_dd\[3\] clknet_leaf_49_clk_regs
+ sg13g2_dfrbpq_1
X_3301_ _1302_ _1301_ _1287_ _1298_ net812 VPWR VGND sg13g2_a22oi_1
X_4281_ net656 VGND VPWR net128 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[43\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
X_3232_ _1243_ VPWR _0233_ VGND _1155_ _1182_ sg13g2_o21ai_1
X_3163_ _1207_ net180 net608 VPWR VGND sg13g2_nand2_1
X_2114_ VPWR _1971_ u_usb_cdc.u_ctrl_endp.in_endp_q VGND sg13g2_inv_1
XFILLER_39_346 VPWR VGND sg13g2_fill_1
X_3094_ _1161_ VPWR _0176_ VGND net828 _1162_ sg13g2_o21ai_1
XFILLER_35_552 VPWR VGND sg13g2_fill_1
XFILLER_35_563 VPWR VGND sg13g2_decap_4
X_3996_ VGND VPWR net904 _1830_ _1831_ net643 sg13g2_a21oi_1
XFILLER_10_419 VPWR VGND sg13g2_decap_8
X_2947_ net509 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ _1077_ _0114_ VPWR VGND sg13g2_mux2_1
X_2878_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net433 _1036_ _0086_ VPWR VGND sg13g2_mux2_1
Xhold420 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[61\] VPWR VGND
+ net463 sg13g2_dlygate4sd3_1
Xhold453 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[7\] VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold442 u_usb_cdc.u_ctrl_endp.addr_dd\[1\] VPWR VGND net485 sg13g2_dlygate4sd3_1
Xhold431 _0280_ VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold475 _0140_ VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold464 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[56\] VPWR VGND
+ net507 sg13g2_dlygate4sd3_1
Xhold486 _0110_ VPWR VGND net529 sg13g2_dlygate4sd3_1
X_4479_ net729 VGND VPWR net267 u_usb_cdc.u_sie.rx_data\[3\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_1
Xhold497 _0336_ VPWR VGND net540 sg13g2_dlygate4sd3_1
XFILLER_26_574 VPWR VGND sg13g2_decap_4
XFILLER_13_213 VPWR VGND sg13g2_fill_2
XFILLER_14_725 VPWR VGND sg13g2_fill_2
XFILLER_26_585 VPWR VGND sg13g2_fill_1
XFILLER_16_1011 VPWR VGND sg13g2_decap_8
XFILLER_10_942 VPWR VGND sg13g2_decap_4
XFILLER_10_997 VPWR VGND sg13g2_decap_8
XFILLER_6_979 VPWR VGND sg13g2_decap_8
XFILLER_0_150 VPWR VGND sg13g2_decap_8
XFILLER_49_611 VPWR VGND sg13g2_decap_8
XFILLER_37_828 VPWR VGND sg13g2_fill_1
XFILLER_49_688 VPWR VGND sg13g2_decap_8
XFILLER_45_883 VPWR VGND sg13g2_decap_8
XFILLER_32_522 VPWR VGND sg13g2_fill_2
X_3850_ _0899_ _1729_ net421 _1732_ VPWR VGND sg13g2_nand3_1
X_2801_ net519 u_usb_cdc.u_sie.data_q\[3\] _2017_ _0854_ _0977_ VPWR VGND sg13g2_nor4_1
XFILLER_32_577 VPWR VGND sg13g2_decap_4
X_3781_ VGND VPWR net810 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[47\]
+ _1680_ _1679_ sg13g2_a21oi_1
XFILLER_9_740 VPWR VGND sg13g2_fill_1
X_2732_ net872 net924 _0925_ VPWR VGND sg13g2_nor2_1
X_2663_ _0864_ _0870_ _0871_ VPWR VGND sg13g2_nor2_1
X_2594_ _0813_ VPWR _0814_ VGND _0650_ _0695_ sg13g2_o21ai_1
X_4402_ net695 VGND VPWR net891 u_usb_cdc.u_sie.crc16_q\[7\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
X_4333_ net681 VGND VPWR _0261_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[2\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_2
X_4264_ net672 VGND VPWR net291 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[26\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_3215_ _1235_ net276 net604 VPWR VGND sg13g2_nand2_1
X_4195_ net666 VGND VPWR net65 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[41\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
X_3146_ net761 net605 _1198_ VPWR VGND sg13g2_nor2_1
XFILLER_39_154 VPWR VGND sg13g2_fill_2
X_3077_ _1149_ net255 net635 VPWR VGND sg13g2_nand2_1
XFILLER_42_319 VPWR VGND sg13g2_decap_8
X_3979_ _1818_ net236 net613 VPWR VGND sg13g2_nand2_1
Xhold261 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[4\] VPWR VGND
+ net304 sg13g2_dlygate4sd3_1
Xhold250 _0414_ VPWR VGND net293 sg13g2_dlygate4sd3_1
XFILLER_49_12 VPWR VGND sg13g2_decap_8
Xhold272 _0032_ VPWR VGND net315 sg13g2_dlygate4sd3_1
Xhold283 _0185_ VPWR VGND net326 sg13g2_dlygate4sd3_1
Xhold294 _0372_ VPWR VGND net337 sg13g2_dlygate4sd3_1
XFILLER_49_89 VPWR VGND sg13g2_fill_1
Xfanout741 net749 net741 VPWR VGND sg13g2_buf_8
Xfanout730 net731 net730 VPWR VGND sg13g2_buf_8
Xfanout763 net764 net763 VPWR VGND sg13g2_buf_8
Xfanout752 net753 net752 VPWR VGND sg13g2_buf_8
Xfanout785 net786 net785 VPWR VGND sg13g2_buf_2
Xfanout774 net775 net774 VPWR VGND sg13g2_buf_1
Xfanout796 net797 net796 VPWR VGND sg13g2_buf_8
XFILLER_46_669 VPWR VGND sg13g2_decap_8
XFILLER_41_352 VPWR VGND sg13g2_fill_1
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_2_982 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_4_clk_regs clknet_3_0__leaf_clk_regs clknet_leaf_4_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3000_ _1111_ VPWR _0133_ VGND _1066_ net610 sg13g2_o21ai_1
Xinput7 ui_in[5] net7 VPWR VGND sg13g2_buf_1
XFILLER_49_485 VPWR VGND sg13g2_decap_8
XFILLER_45_691 VPWR VGND sg13g2_decap_8
X_3902_ net457 _1765_ _1769_ VPWR VGND sg13g2_and2_1
X_3833_ VPWR _1719_ _1718_ VGND sg13g2_inv_1
X_3764_ _1663_ VPWR _1664_ VGND net807 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[38\]
+ sg13g2_o21ai_1
X_2715_ net990 _2043_ _0429_ _0913_ VPWR VGND sg13g2_nor3_1
X_3695_ _1591_ VPWR _1598_ VGND _1594_ _1597_ sg13g2_o21ai_1
X_2646_ _0857_ net710 _0856_ VPWR VGND sg13g2_nand2_1
X_2577_ _0694_ _0706_ _0802_ VPWR VGND u_usb_cdc.u_ctrl_endp.in_dir_q sg13g2_nand3b_1
X_4316_ net648 VGND VPWR net260 net21 clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
X_4247_ net658 VGND VPWR net104 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[9\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_4178_ net680 VGND VPWR net516 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[24\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
X_3129_ VGND VPWR net632 _1186_ _0187_ _1185_ sg13g2_a21oi_1
XFILLER_27_168 VPWR VGND sg13g2_decap_8
XFILLER_28_669 VPWR VGND sg13g2_fill_1
XFILLER_42_105 VPWR VGND sg13g2_fill_2
XFILLER_13_1003 VPWR VGND sg13g2_decap_8
XFILLER_3_724 VPWR VGND sg13g2_decap_8
XFILLER_47_901 VPWR VGND sg13g2_decap_8
Xfanout582 _1401_ net582 VPWR VGND sg13g2_buf_1
Xfanout593 net594 net593 VPWR VGND sg13g2_buf_8
XFILLER_18_102 VPWR VGND sg13g2_fill_1
XFILLER_19_658 VPWR VGND sg13g2_decap_8
XFILLER_20_1018 VPWR VGND sg13g2_decap_8
XFILLER_47_978 VPWR VGND sg13g2_decap_8
XFILLER_27_680 VPWR VGND sg13g2_fill_1
XFILLER_33_149 VPWR VGND sg13g2_fill_2
XFILLER_15_886 VPWR VGND sg13g2_decap_4
XFILLER_42_661 VPWR VGND sg13g2_fill_1
XFILLER_41_193 VPWR VGND sg13g2_fill_2
X_2500_ _0727_ net723 u_usb_cdc.sie_out_data\[1\] VPWR VGND sg13g2_nand2_1
X_3480_ u_usb_cdc.sie_out_data\[5\] _1421_ _1432_ VPWR VGND sg13g2_nor2_1
X_2431_ _0661_ _0633_ _0660_ VPWR VGND sg13g2_nand2_2
X_2362_ u_usb_cdc.sie_in_data_ack u_usb_cdc.sie_in_req _0593_ VPWR VGND sg13g2_nor2_1
X_4101_ net686 VGND VPWR net958 u_usb_cdc.u_ctrl_endp.req_q\[7\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_2
X_2293_ net787 u_usb_cdc.u_ctrl_endp.max_length_q\[2\] _0525_ VPWR VGND sg13g2_xor2_1
X_4032_ VPWR VGND _1823_ _1822_ _1862_ u_usb_cdc.u_sie.u_phy_tx.data_q\[5\] _1863_
+ _1830_ sg13g2_a221oi_1
XFILLER_38_945 VPWR VGND sg13g2_decap_8
XFILLER_49_293 VPWR VGND sg13g2_decap_4
XFILLER_49_282 VPWR VGND sg13g2_fill_2
XFILLER_36_1014 VPWR VGND sg13g2_decap_8
X_3816_ _0862_ _1701_ net488 _1706_ VPWR VGND sg13g2_nand3_1
X_3747_ net800 VPWR _1648_ VGND net805 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[53\]
+ sg13g2_o21ai_1
X_3678_ _1574_ VPWR _1582_ VGND net795 _1581_ sg13g2_o21ai_1
X_2629_ VGND VPWR _0841_ _0481_ _0453_ sg13g2_or2_1
XFILLER_0_727 VPWR VGND sg13g2_decap_8
XFILLER_29_945 VPWR VGND sg13g2_decap_8
XFILLER_16_606 VPWR VGND sg13g2_fill_1
XFILLER_46_68 VPWR VGND sg13g2_fill_1
XFILLER_11_377 VPWR VGND sg13g2_decap_4
XFILLER_3_554 VPWR VGND sg13g2_decap_8
XFILLER_4_1023 VPWR VGND sg13g2_decap_4
XFILLER_47_775 VPWR VGND sg13g2_decap_8
X_2980_ _1101_ net64 _1096_ VPWR VGND sg13g2_nand2_1
XFILLER_30_642 VPWR VGND sg13g2_decap_8
X_3601_ _1507_ _0539_ _0670_ VPWR VGND sg13g2_nand2_1
Xinput10 uio_in[0] net10 VPWR VGND sg13g2_buf_1
X_3532_ VGND VPWR _1917_ net585 _0312_ _1464_ sg13g2_a21oi_1
XFILLER_7_893 VPWR VGND sg13g2_fill_1
X_3463_ net881 net576 _1420_ VPWR VGND sg13g2_nor2_1
X_2414_ VPWR _0644_ _0643_ VGND sg13g2_inv_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
X_3394_ net419 _1133_ _1378_ VPWR VGND sg13g2_nor2_1
X_2345_ VGND VPWR _0482_ _0576_ _0577_ net752 sg13g2_a21oi_1
XFILLER_29_208 VPWR VGND sg13g2_fill_2
X_2276_ _0502_ _0503_ _0496_ _0508_ VPWR VGND _0504_ sg13g2_nand4_1
X_4015_ _2028_ _1846_ _1847_ _1848_ VPWR VGND sg13g2_nor3_1
XFILLER_37_252 VPWR VGND sg13g2_fill_1
XFILLER_16_49 VPWR VGND sg13g2_fill_1
XFILLER_12_119 VPWR VGND sg13g2_fill_1
XFILLER_0_568 VPWR VGND sg13g2_decap_8
XFILLER_48_506 VPWR VGND sg13g2_decap_8
XFILLER_29_786 VPWR VGND sg13g2_fill_2
XFILLER_44_767 VPWR VGND sg13g2_decap_8
XFILLER_32_918 VPWR VGND sg13g2_decap_8
XFILLER_24_491 VPWR VGND sg13g2_fill_1
Xheichips25_usb_cdc_33 VPWR VGND uio_oe[1] sg13g2_tielo
XFILLER_26_1002 VPWR VGND sg13g2_decap_8
X_2130_ VPWR _0039_ net49 VGND sg13g2_inv_1
X_2061_ VPWR _1918_ net1037 VGND sg13g2_inv_1
X_2963_ _1089_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net636 VPWR VGND sg13g2_nand2_1
XFILLER_15_491 VPWR VGND sg13g2_decap_8
X_2894_ _1045_ VPWR _0092_ VGND net618 _1046_ sg13g2_o21ai_1
XFILLER_31_995 VPWR VGND sg13g2_decap_8
Xhold602 u_usb_cdc.u_sie.phy_state_q\[6\] VPWR VGND net921 sg13g2_dlygate4sd3_1
Xhold635 _0285_ VPWR VGND net954 sg13g2_dlygate4sd3_1
Xhold613 u_usb_cdc.u_sie.crc16_q\[1\] VPWR VGND net932 sg13g2_dlygate4sd3_1
X_3515_ _1264_ _1457_ _0302_ VPWR VGND sg13g2_and2_1
Xhold624 _0004_ VPWR VGND net943 sg13g2_dlygate4sd3_1
Xhold646 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[3\] VPWR
+ VGND net965 sg13g2_dlygate4sd3_1
Xhold668 _0580_ VPWR VGND net987 sg13g2_dlygate4sd3_1
Xhold679 u_usb_cdc.u_sie.pid_q\[2\] VPWR VGND net998 sg13g2_dlygate4sd3_1
X_4495_ net701 VGND VPWR _0412_ u_usb_cdc.u_sie.u_phy_tx.data_q\[2\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
Xhold657 u_usb_cdc.u_sie.u_phy_rx.rx_en_q VPWR VGND net976 sg13g2_dlygate4sd3_1
X_3446_ _1940_ _0640_ _0693_ _1409_ VPWR VGND sg13g2_nor3_1
X_3377_ _0257_ net813 _1363_ VPWR VGND sg13g2_xnor2_1
X_2328_ _0560_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[1\] net801
+ VPWR VGND sg13g2_xnor2_1
XFILLER_45_509 VPWR VGND sg13g2_decap_4
X_2259_ _0491_ u_usb_cdc.u_sie.crc16_q\[13\] net765 VPWR VGND sg13g2_xnor2_1
XFILLER_38_583 VPWR VGND sg13g2_decap_8
XFILLER_43_47 VPWR VGND sg13g2_fill_1
XFILLER_43_69 VPWR VGND sg13g2_fill_1
XFILLER_49_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_19 VPWR VGND sg13g2_fill_1
XFILLER_1_811 VPWR VGND sg13g2_decap_8
XFILLER_0_365 VPWR VGND sg13g2_decap_8
XFILLER_17_701 VPWR VGND sg13g2_fill_2
XFILLER_29_594 VPWR VGND sg13g2_decap_8
XFILLER_31_236 VPWR VGND sg13g2_fill_2
XFILLER_9_922 VPWR VGND sg13g2_decap_4
XFILLER_9_988 VPWR VGND sg13g2_decap_8
X_3300_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[1\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[9\]
+ net824 _1301_ VPWR VGND sg13g2_mux2_1
X_4280_ net654 VGND VPWR net176 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[42\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_3231_ _1243_ net207 _1156_ VPWR VGND sg13g2_nand2_1
X_3162_ _1206_ VPWR _0200_ VGND _1180_ net609 sg13g2_o21ai_1
X_2113_ VPWR _1970_ net418 VGND sg13g2_inv_1
XFILLER_12_2 VPWR VGND sg13g2_fill_1
X_3093_ net832 _1159_ net762 _1162_ VPWR VGND sg13g2_nand3_1
XFILLER_48_892 VPWR VGND sg13g2_decap_8
X_3995_ _2020_ _1008_ _1830_ VPWR VGND sg13g2_and2_1
X_2946_ net570 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ _1077_ _0113_ VPWR VGND sg13g2_mux2_1
X_2877_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net490 _1036_ _0085_ VPWR VGND sg13g2_mux2_1
Xhold410 _1811_ VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold443 u_usb_cdc.u_sie.out_toggle_q\[0\] VPWR VGND net486 sg13g2_dlygate4sd3_1
Xhold432 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[60\] VPWR VGND
+ net475 sg13g2_dlygate4sd3_1
Xhold421 _0144_ VPWR VGND net464 sg13g2_dlygate4sd3_1
Xhold454 _0367_ VPWR VGND net497 sg13g2_dlygate4sd3_1
Xhold487 u_usb_cdc.u_sie.crc16_q\[0\] VPWR VGND net530 sg13g2_dlygate4sd3_1
Xhold465 _0139_ VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold476 u_usb_cdc.u_sie.data_q\[2\] VPWR VGND net519 sg13g2_dlygate4sd3_1
X_4478_ net729 VGND VPWR net233 u_usb_cdc.u_sie.rx_data\[2\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_1
X_3429_ u_usb_cdc.sie_out_data\[7\] _1941_ _0640_ _1399_ VPWR VGND sg13g2_nor3_1
Xhold498 _0049_ VPWR VGND net541 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_28_clk_regs clknet_3_7__leaf_clk_regs clknet_leaf_28_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_45_317 VPWR VGND sg13g2_decap_4
XFILLER_14_704 VPWR VGND sg13g2_decap_8
XFILLER_13_269 VPWR VGND sg13g2_fill_2
XFILLER_22_781 VPWR VGND sg13g2_fill_2
XFILLER_6_914 VPWR VGND sg13g2_fill_1
XFILLER_5_435 VPWR VGND sg13g2_fill_2
XFILLER_6_958 VPWR VGND sg13g2_decap_8
XFILLER_1_685 VPWR VGND sg13g2_decap_8
XFILLER_23_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_667 VPWR VGND sg13g2_decap_8
XFILLER_45_862 VPWR VGND sg13g2_decap_8
X_2800_ _0975_ VPWR _0976_ VGND net839 net844 sg13g2_o21ai_1
XFILLER_32_589 VPWR VGND sg13g2_fill_1
X_3780_ net810 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[39\] _1679_
+ VPWR VGND sg13g2_nor2b_1
X_2731_ net626 _0923_ _0924_ VPWR VGND sg13g2_nor2_1
XFILLER_8_284 VPWR VGND sg13g2_fill_2
X_2662_ net844 VPWR _0870_ VGND u_usb_cdc.u_sie.data_q\[1\] _0863_ sg13g2_o21ai_1
X_4401_ net700 VGND VPWR net907 u_usb_cdc.u_sie.crc16_q\[6\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
X_2593_ _0813_ _0673_ _0692_ VPWR VGND sg13g2_nand2_1
XFILLER_5_991 VPWR VGND sg13g2_decap_8
X_4332_ net681 VGND VPWR net1016 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[1\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_1
X_4263_ net672 VGND VPWR _0192_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[25\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_3214_ net101 VPWR _0224_ VGND net722 net604 sg13g2_o21ai_1
X_4194_ net680 VGND VPWR net63 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[40\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
X_3145_ _1197_ VPWR _0192_ VGND net722 net606 sg13g2_o21ai_1
X_3076_ _1148_ VPWR _0172_ VGND _1914_ net634 sg13g2_o21ai_1
XFILLER_39_1023 VPWR VGND sg13g2_decap_4
XFILLER_11_718 VPWR VGND sg13g2_decap_8
X_3978_ _1817_ VPWR _0405_ VGND _1950_ net613 sg13g2_o21ai_1
X_2929_ _1069_ VPWR _0103_ VGND net619 _1070_ sg13g2_o21ai_1
Xhold262 u_usb_cdc.u_sie.u_phy_rx.rx_err_q VPWR VGND net305 sg13g2_dlygate4sd3_1
Xhold251 net25 VPWR VGND net294 sg13g2_dlygate4sd3_1
Xhold240 _0376_ VPWR VGND net283 sg13g2_dlygate4sd3_1
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_1016 VPWR VGND sg13g2_decap_8
Xhold273 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[20\] VPWR
+ VGND net316 sg13g2_dlygate4sd3_1
Xhold284 u_usb_cdc.u_sie.in_byte_q\[0\] VPWR VGND net327 sg13g2_dlygate4sd3_1
Xhold295 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[6\] VPWR VGND net338 sg13g2_dlygate4sd3_1
Xfanout720 _1912_ net720 VPWR VGND sg13g2_buf_8
Xfanout742 net743 net742 VPWR VGND sg13g2_buf_8
XFILLER_49_68 VPWR VGND sg13g2_decap_8
Xfanout731 net732 net731 VPWR VGND sg13g2_buf_8
Xfanout764 u_usb_cdc.sie_out_data\[0\] net764 VPWR VGND sg13g2_buf_8
Xfanout753 net754 net753 VPWR VGND sg13g2_buf_8
Xfanout775 net1049 net775 VPWR VGND sg13g2_buf_8
Xfanout786 net787 net786 VPWR VGND sg13g2_buf_1
Xfanout797 net1040 net797 VPWR VGND sg13g2_buf_8
XFILLER_46_648 VPWR VGND sg13g2_decap_8
XFILLER_45_169 VPWR VGND sg13g2_fill_2
XFILLER_14_512 VPWR VGND sg13g2_fill_1
XFILLER_27_895 VPWR VGND sg13g2_decap_8
XFILLER_6_700 VPWR VGND sg13g2_decap_8
XFILLER_5_254 VPWR VGND sg13g2_fill_2
XFILLER_2_961 VPWR VGND sg13g2_decap_8
XFILLER_7_1021 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[6] net8 VPWR VGND sg13g2_buf_1
XFILLER_49_464 VPWR VGND sg13g2_decap_8
XFILLER_33_843 VPWR VGND sg13g2_fill_2
X_3901_ _1768_ net713 net457 VPWR VGND sg13g2_nand2_1
X_3832_ net717 _1717_ _1718_ VPWR VGND sg13g2_nor2_1
X_3763_ VGND VPWR net808 _1991_ _1663_ net800 sg13g2_a21oi_1
X_2714_ VGND VPWR _0912_ _2044_ _2039_ sg13g2_or2_1
X_3694_ net796 VPWR _1597_ VGND _1595_ _1596_ sg13g2_o21ai_1
X_2645_ net765 _0454_ _0855_ _0856_ VPWR VGND sg13g2_nor3_1
X_2576_ net483 VPWR _0801_ VGND _0795_ _0800_ sg13g2_o21ai_1
X_4315_ net648 VGND VPWR net297 net20 clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
XFILLER_0_909 VPWR VGND sg13g2_decap_8
XFILLER_19_38 VPWR VGND sg13g2_fill_1
X_4246_ net658 VGND VPWR net204 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[8\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_4177_ net669 VGND VPWR net122 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[23\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_3128_ _1186_ net759 _1141_ VPWR VGND sg13g2_nand2_2
X_3059_ _1138_ net363 _1135_ VPWR VGND sg13g2_nand2_1
XFILLER_24_843 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_43_clk_regs clknet_3_4__leaf_clk_regs clknet_leaf_43_clk_regs VPWR VGND
+ sg13g2_buf_8
Xfanout583 net584 net583 VPWR VGND sg13g2_buf_8
XFILLER_47_957 VPWR VGND sg13g2_decap_8
Xfanout594 _0521_ net594 VPWR VGND sg13g2_buf_8
XFILLER_34_607 VPWR VGND sg13g2_fill_1
XFILLER_33_117 VPWR VGND sg13g2_fill_1
XFILLER_6_585 VPWR VGND sg13g2_decap_4
X_2430_ _0654_ _0658_ _0659_ _0660_ VPWR VGND sg13g2_nor3_1
XFILLER_29_1022 VPWR VGND sg13g2_decap_8
X_2361_ _0435_ VPWR _0592_ VGND _0587_ _0591_ sg13g2_o21ai_1
X_4100_ net689 VGND VPWR net484 u_usb_cdc.u_ctrl_endp.req_q\[6\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_2
X_2292_ net779 u_usb_cdc.u_ctrl_endp.max_length_q\[3\] _0524_ VPWR VGND sg13g2_xor2_1
XFILLER_1_290 VPWR VGND sg13g2_decap_8
X_4031_ _1860_ _1861_ _1859_ _1862_ VPWR VGND sg13g2_nand3_1
X_3815_ _1705_ net848 _1704_ VPWR VGND sg13g2_nand2_1
X_3746_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[61\] net805 _1647_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_21_39 VPWR VGND sg13g2_decap_8
X_3677_ _1580_ VPWR _1581_ VGND net796 _1575_ sg13g2_o21ai_1
X_2628_ _0840_ net847 net596 VPWR VGND sg13g2_nand2_1
XFILLER_0_706 VPWR VGND sg13g2_decap_8
X_2559_ _0757_ _0785_ _0721_ _0004_ VPWR VGND sg13g2_nand3_1
X_4229_ net661 VGND VPWR _0158_ u_usb_cdc.in_ready_o[0] clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
XFILLER_29_924 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_46_47 VPWR VGND sg13g2_fill_1
XFILLER_44_949 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_fill_1
XFILLER_30_109 VPWR VGND sg13g2_fill_2
XFILLER_23_172 VPWR VGND sg13g2_fill_1
XFILLER_24_684 VPWR VGND sg13g2_decap_8
XFILLER_7_316 VPWR VGND sg13g2_fill_2
XFILLER_4_1002 VPWR VGND sg13g2_decap_8
XFILLER_35_905 VPWR VGND sg13g2_fill_1
XFILLER_47_754 VPWR VGND sg13g2_decap_8
XFILLER_43_982 VPWR VGND sg13g2_decap_8
XFILLER_15_640 VPWR VGND sg13g2_fill_2
XFILLER_21_109 VPWR VGND sg13g2_fill_1
X_3600_ _1506_ net780 _0539_ VPWR VGND sg13g2_nand2_2
XFILLER_30_698 VPWR VGND sg13g2_fill_1
Xinput11 uio_in[1] net11 VPWR VGND sg13g2_buf_1
X_3531_ net409 net585 _1464_ VPWR VGND sg13g2_nor2_1
XFILLER_6_382 VPWR VGND sg13g2_fill_2
X_3462_ _1389_ _1418_ _1419_ VPWR VGND sg13g2_nor2_1
X_2413_ net849 u_usb_cdc.u_ctrl_endp.state_q\[6\] _0551_ _0643_ VPWR VGND sg13g2_nor3_1
X_3393_ net1015 VPWR _0260_ VGND _1369_ _1376_ sg13g2_o21ai_1
X_2344_ _0513_ _0575_ _0576_ VPWR VGND sg13g2_and2_1
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk VPWR VGND sg13g2_buf_8
X_2275_ _0500_ _0505_ _0499_ _0507_ VPWR VGND sg13g2_nand3_1
X_4014_ _1842_ VPWR _1847_ VGND net383 _1835_ sg13g2_o21ai_1
XFILLER_26_938 VPWR VGND sg13g2_fill_2
XFILLER_37_275 VPWR VGND sg13g2_fill_1
XFILLER_40_429 VPWR VGND sg13g2_fill_2
XFILLER_20_131 VPWR VGND sg13g2_fill_2
XFILLER_32_16 VPWR VGND sg13g2_decap_8
XFILLER_21_698 VPWR VGND sg13g2_fill_2
XFILLER_4_319 VPWR VGND sg13g2_fill_1
XFILLER_10_1018 VPWR VGND sg13g2_decap_8
X_3729_ _1627_ _1628_ _1631_ VPWR VGND _1629_ sg13g2_nand3b_1
XFILLER_0_547 VPWR VGND sg13g2_decap_8
XFILLER_28_242 VPWR VGND sg13g2_fill_1
XFILLER_28_253 VPWR VGND sg13g2_fill_2
XFILLER_44_746 VPWR VGND sg13g2_decap_8
XFILLER_43_278 VPWR VGND sg13g2_decap_4
XFILLER_8_603 VPWR VGND sg13g2_decap_8
XFILLER_40_985 VPWR VGND sg13g2_decap_8
XFILLER_8_647 VPWR VGND sg13g2_decap_4
XFILLER_4_820 VPWR VGND sg13g2_decap_4
Xheichips25_usb_cdc_34 VPWR VGND uio_oe[2] sg13g2_tielo
X_2060_ net758 _1917_ VPWR VGND sg13g2_inv_4
X_2962_ _1088_ net205 _1079_ VPWR VGND sg13g2_nand2_1
X_2893_ _1046_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net645 VPWR VGND sg13g2_nand2_1
XFILLER_31_974 VPWR VGND sg13g2_decap_8
XFILLER_30_484 VPWR VGND sg13g2_decap_4
Xhold603 u_usb_cdc.u_ctrl_endp.max_length_q\[4\] VPWR VGND net922 sg13g2_dlygate4sd3_1
Xhold636 u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] VPWR VGND net955 sg13g2_dlygate4sd3_1
Xhold625 u_usb_cdc.u_sie.pid_q\[1\] VPWR VGND net944 sg13g2_dlygate4sd3_1
X_4494_ net702 VGND VPWR _0411_ u_usb_cdc.u_sie.u_phy_tx.data_q\[1\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
X_3514_ _1457_ _1249_ net770 VPWR VGND sg13g2_nand2b_1
Xhold614 u_usb_cdc.in_ready_o[0] VPWR VGND net933 sg13g2_dlygate4sd3_1
X_3445_ VGND VPWR _1917_ net581 _0281_ _1408_ sg13g2_a21oi_1
Xhold669 _0581_ VPWR VGND net988 sg13g2_dlygate4sd3_1
Xhold647 _0258_ VPWR VGND net966 sg13g2_dlygate4sd3_1
Xhold658 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[0\] VPWR VGND
+ net977 sg13g2_dlygate4sd3_1
X_3376_ _1363_ _1364_ _0256_ VPWR VGND sg13g2_and2_1
X_2327_ _0559_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[2\] net797
+ VPWR VGND sg13g2_xnor2_1
X_2258_ _0490_ _0485_ _0488_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_49 VPWR VGND sg13g2_decap_8
X_2189_ _2043_ net976 _2040_ VPWR VGND sg13g2_nand2_1
XFILLER_26_735 VPWR VGND sg13g2_fill_1
XFILLER_14_908 VPWR VGND sg13g2_fill_1
XFILLER_21_484 VPWR VGND sg13g2_decap_4
XFILLER_49_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_344 VPWR VGND sg13g2_decap_8
XFILLER_49_849 VPWR VGND sg13g2_decap_8
XFILLER_17_71 VPWR VGND sg13g2_decap_4
XFILLER_13_963 VPWR VGND sg13g2_fill_2
XFILLER_13_952 VPWR VGND sg13g2_fill_1
XFILLER_12_440 VPWR VGND sg13g2_fill_1
XFILLER_13_996 VPWR VGND sg13g2_decap_8
XFILLER_9_967 VPWR VGND sg13g2_decap_8
XFILLER_8_488 VPWR VGND sg13g2_decap_4
XFILLER_3_160 VPWR VGND sg13g2_fill_2
X_3230_ _1242_ VPWR _0232_ VGND _1155_ _1180_ sg13g2_o21ai_1
X_3161_ _1206_ net143 net609 VPWR VGND sg13g2_nand2_1
X_2112_ _1969_ net906 VPWR VGND sg13g2_inv_2
XFILLER_48_871 VPWR VGND sg13g2_decap_8
X_3092_ _1161_ net103 _1151_ VPWR VGND sg13g2_nand2_1
XFILLER_35_543 VPWR VGND sg13g2_fill_2
XFILLER_23_716 VPWR VGND sg13g2_decap_8
X_3994_ _1008_ _1827_ _1828_ _1829_ VPWR VGND sg13g2_or3_1
X_2945_ net520 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ _1077_ _0112_ VPWR VGND sg13g2_mux2_1
X_2876_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net549 _1036_ _0084_ VPWR VGND sg13g2_mux2_1
Xhold411 _0398_ VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold400 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[4\] VPWR VGND
+ net443 sg13g2_dlygate4sd3_1
Xhold444 _0067_ VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold422 u_usb_cdc.u_sie.u_phy_rx.rx_eop_qq VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold433 _0143_ VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold455 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[52\] VPWR
+ VGND net498 sg13g2_dlygate4sd3_1
X_4477_ net730 VGND VPWR _0402_ u_usb_cdc.u_sie.rx_data\[1\] clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_1
Xhold477 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[29\] VPWR VGND
+ net520 sg13g2_dlygate4sd3_1
Xhold466 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[31\] VPWR VGND
+ net509 sg13g2_dlygate4sd3_1
Xhold488 _0323_ VPWR VGND net531 sg13g2_dlygate4sd3_1
X_3428_ VGND VPWR net850 _0601_ _1398_ net715 sg13g2_a21oi_1
Xhold499 _0062_ VPWR VGND net542 sg13g2_dlygate4sd3_1
X_3359_ _1353_ VPWR _1354_ VGND net824 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[7\]
+ sg13g2_o21ai_1
XFILLER_38_15 VPWR VGND sg13g2_fill_2
XFILLER_38_48 VPWR VGND sg13g2_fill_2
XFILLER_41_557 VPWR VGND sg13g2_decap_4
XFILLER_10_922 VPWR VGND sg13g2_decap_8
XFILLER_1_664 VPWR VGND sg13g2_decap_8
XFILLER_23_1006 VPWR VGND sg13g2_decap_8
XFILLER_49_646 VPWR VGND sg13g2_decap_8
XFILLER_48_167 VPWR VGND sg13g2_fill_1
XFILLER_45_841 VPWR VGND sg13g2_decap_8
XFILLER_17_587 VPWR VGND sg13g2_fill_2
XFILLER_32_524 VPWR VGND sg13g2_fill_1
XFILLER_32_546 VPWR VGND sg13g2_fill_2
XFILLER_9_731 VPWR VGND sg13g2_decap_4
X_2730_ _0923_ net625 net709 VPWR VGND sg13g2_nand2_2
X_2661_ _0869_ VPWR _0023_ VGND _0587_ _0867_ sg13g2_o21ai_1
X_4400_ net700 VGND VPWR _0328_ u_usb_cdc.u_sie.crc16_q\[5\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
X_2592_ _0794_ _0796_ _0701_ _0812_ VPWR VGND _0799_ sg13g2_nand4_1
XFILLER_5_970 VPWR VGND sg13g2_decap_8
X_4331_ net681 VGND VPWR _0259_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[0\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_1
X_4262_ net672 VGND VPWR net173 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[24\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_3213_ _1234_ net100 _1232_ VPWR VGND sg13g2_nand2_1
X_4193_ net669 VGND VPWR net178 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[39\]
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
X_3144_ _1197_ net145 net606 VPWR VGND sg13g2_nand2_1
XFILLER_10_0 VPWR VGND sg13g2_fill_2
XFILLER_39_156 VPWR VGND sg13g2_fill_1
X_3075_ _1148_ net286 net634 VPWR VGND sg13g2_nand2_1
XFILLER_39_1002 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_fill_2
X_3977_ _1817_ net228 net613 VPWR VGND sg13g2_nand2_1
X_2928_ _1070_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net644 VPWR VGND sg13g2_nand2_1
X_2859_ _1026_ _1027_ _1024_ _1030_ VPWR VGND _1029_ sg13g2_nand4_1
XFILLER_3_918 VPWR VGND sg13g2_fill_2
Xhold230 _0196_ VPWR VGND net273 sg13g2_dlygate4sd3_1
Xhold252 _0249_ VPWR VGND net295 sg13g2_dlygate4sd3_1
X_4529_ u_usb_cdc.out_valid_o[0] net15 VPWR VGND sg13g2_buf_1
Xhold241 u_usb_cdc.u_sie.rx_data\[1\] VPWR VGND net284 sg13g2_dlygate4sd3_1
Xhold263 _0944_ VPWR VGND net306 sg13g2_dlygate4sd3_1
Xhold274 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[48\] VPWR
+ VGND net317 sg13g2_dlygate4sd3_1
Xhold285 _0319_ VPWR VGND net328 sg13g2_dlygate4sd3_1
Xhold296 _0366_ VPWR VGND net339 sg13g2_dlygate4sd3_1
Xfanout732 net738 net732 VPWR VGND sg13g2_buf_8
Xfanout721 net722 net721 VPWR VGND sg13g2_buf_8
Xfanout710 _2015_ net710 VPWR VGND sg13g2_buf_8
XFILLER_49_47 VPWR VGND sg13g2_decap_8
Xfanout765 net519 net765 VPWR VGND sg13g2_buf_8
Xfanout743 net744 net743 VPWR VGND sg13g2_buf_8
Xfanout754 net876 net754 VPWR VGND sg13g2_buf_8
Xfanout776 net778 net776 VPWR VGND sg13g2_buf_8
Xfanout798 net800 net798 VPWR VGND sg13g2_buf_8
Xfanout787 net1050 net787 VPWR VGND sg13g2_buf_8
XFILLER_27_830 VPWR VGND sg13g2_decap_4
XFILLER_6_745 VPWR VGND sg13g2_fill_2
XFILLER_2_940 VPWR VGND sg13g2_decap_8
XFILLER_1_461 VPWR VGND sg13g2_decap_8
XFILLER_7_1000 VPWR VGND sg13g2_decap_8
XFILLER_49_443 VPWR VGND sg13g2_decap_8
Xinput9 ui_in[7] net9 VPWR VGND sg13g2_buf_1
XFILLER_37_627 VPWR VGND sg13g2_fill_2
X_3900_ net879 net713 _1767_ _0377_ VPWR VGND sg13g2_a21o_1
X_3831_ _0436_ _0603_ _1474_ _1717_ VPWR VGND sg13g2_mux2_1
X_3762_ net804 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[6\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[14\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[22\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[30\]
+ net798 _1662_ VPWR VGND sg13g2_mux4_1
X_2713_ _0905_ _0908_ _0902_ _0030_ VPWR VGND _0911_ sg13g2_nand4_1
X_3693_ net799 VPWR _1596_ VGND net803 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[51\]
+ sg13g2_o21ai_1
X_2644_ _0451_ VPWR _0855_ VGND u_usb_cdc.u_sie.pid_q\[2\] _1935_ sg13g2_o21ai_1
X_2575_ _0797_ _0798_ _0796_ _0800_ VPWR VGND _0799_ sg13g2_nand4_1
X_4314_ net648 VGND VPWR _0243_ net19 clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
X_4245_ net658 VGND VPWR _0174_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[7\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_4176_ net670 VGND VPWR net239 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[22\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_3127_ net316 net632 _1185_ VPWR VGND sg13g2_nor2_1
XFILLER_42_107 VPWR VGND sg13g2_fill_1
XFILLER_42_118 VPWR VGND sg13g2_fill_2
X_3058_ _1137_ VPWR _0165_ VGND _1923_ _1135_ sg13g2_o21ai_1
XFILLER_36_660 VPWR VGND sg13g2_fill_2
Xfanout584 _1492_ net584 VPWR VGND sg13g2_buf_8
XFILLER_47_936 VPWR VGND sg13g2_decap_8
Xfanout595 _0901_ net595 VPWR VGND sg13g2_buf_8
XFILLER_19_638 VPWR VGND sg13g2_decap_8
XFILLER_46_402 VPWR VGND sg13g2_fill_2
XFILLER_18_126 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_12_clk_regs clknet_3_3__leaf_clk_regs clknet_leaf_12_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_25_60 VPWR VGND sg13g2_decap_8
Xi_spad_env_f_bit VGND VPWR clknet_1_0__leaf_clk net18 net14 uio_in[2] spad_env_f_bit
XFILLER_6_553 VPWR VGND sg13g2_fill_2
XFILLER_6_564 VPWR VGND sg13g2_fill_1
XFILLER_29_1001 VPWR VGND sg13g2_decap_8
X_2360_ _0556_ _0564_ _0569_ _0589_ _0591_ VPWR VGND sg13g2_nor4_1
X_2291_ _0523_ net844 _0522_ VPWR VGND sg13g2_nand2_1
X_4030_ _1861_ _1964_ net837 u_usb_cdc.u_sie.data_q\[4\] net842 VPWR VGND sg13g2_a22oi_1
XFILLER_2_97 VPWR VGND sg13g2_fill_2
XFILLER_18_693 VPWR VGND sg13g2_decap_4
XFILLER_33_630 VPWR VGND sg13g2_fill_1
XFILLER_33_652 VPWR VGND sg13g2_decap_8
XFILLER_21_814 VPWR VGND sg13g2_decap_8
X_3814_ VGND VPWR u_usb_cdc.ctrl_stall net641 _1704_ _0568_ sg13g2_a21oi_1
X_3745_ net798 _1644_ _1645_ _1646_ VPWR VGND sg13g2_nor3_1
X_3676_ _1580_ _1577_ _1579_ VPWR VGND sg13g2_nand2_1
X_2627_ _0839_ VPWR _0017_ VGND _1928_ _0619_ sg13g2_o21ai_1
X_2558_ _0785_ _0784_ _0662_ _0760_ _0758_ VPWR VGND sg13g2_a22oi_1
X_2489_ net938 _0716_ _0717_ VPWR VGND sg13g2_nor2_2
X_4228_ net681 VGND VPWR net883 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\]
+ clknet_leaf_20_clk_regs sg13g2_dfrbpq_1
X_4159_ net663 VGND VPWR net456 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[5\]
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
XFILLER_44_928 VPWR VGND sg13g2_decap_8
XFILLER_47_733 VPWR VGND sg13g2_decap_8
XFILLER_46_276 VPWR VGND sg13g2_fill_2
XFILLER_43_961 VPWR VGND sg13g2_decap_8
Xinput12 usb_dn_rx_i net12 VPWR VGND sg13g2_buf_1
X_3530_ VGND VPWR _1914_ net586 _0311_ _1463_ sg13g2_a21oi_1
XFILLER_7_840 VPWR VGND sg13g2_fill_1
X_3461_ net624 _0648_ _1417_ _1418_ VPWR VGND sg13g2_nor3_1
X_2412_ _0637_ _0641_ _0642_ VPWR VGND sg13g2_nor2_1
X_3392_ _1377_ net802 _1369_ VPWR VGND sg13g2_nand2_1
X_2343_ VGND VPWR net847 _2017_ _0575_ _0520_ sg13g2_a21oi_1
X_4013_ VGND VPWR _0926_ _1845_ _1846_ _1834_ sg13g2_a21oi_1
X_2274_ _0506_ net840 net751 VPWR VGND sg13g2_nand2b_1
XFILLER_37_210 VPWR VGND sg13g2_fill_2
XFILLER_19_991 VPWR VGND sg13g2_fill_2
XFILLER_21_622 VPWR VGND sg13g2_fill_2
XFILLER_34_994 VPWR VGND sg13g2_decap_8
XFILLER_21_644 VPWR VGND sg13g2_fill_1
XFILLER_21_688 VPWR VGND sg13g2_fill_2
X_3728_ _1630_ _1512_ _1628_ VPWR VGND sg13g2_nand2_1
X_3659_ _1536_ VPWR _0340_ VGND _1562_ _1563_ sg13g2_o21ai_1
XFILLER_0_526 VPWR VGND sg13g2_decap_8
XFILLER_28_210 VPWR VGND sg13g2_fill_1
XFILLER_29_788 VPWR VGND sg13g2_fill_1
XFILLER_44_714 VPWR VGND sg13g2_fill_2
XFILLER_19_1011 VPWR VGND sg13g2_decap_8
XFILLER_12_622 VPWR VGND sg13g2_fill_2
XFILLER_25_983 VPWR VGND sg13g2_decap_8
XFILLER_40_964 VPWR VGND sg13g2_decap_8
XFILLER_22_61 VPWR VGND sg13g2_fill_1
XFILLER_7_158 VPWR VGND sg13g2_fill_1
Xheichips25_usb_cdc_35 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_3_386 VPWR VGND sg13g2_decap_8
XFILLER_16_961 VPWR VGND sg13g2_fill_2
XFILLER_35_758 VPWR VGND sg13g2_fill_1
XFILLER_16_983 VPWR VGND sg13g2_fill_1
X_2961_ _1086_ VPWR _0118_ VGND net618 _1087_ sg13g2_o21ai_1
X_2892_ _1045_ net193 _1037_ VPWR VGND sg13g2_nand2_1
XFILLER_33_1019 VPWR VGND sg13g2_decap_4
Xhold604 u_usb_cdc.addr\[3\] VPWR VGND net923 sg13g2_dlygate4sd3_1
Xhold626 _0356_ VPWR VGND net945 sg13g2_dlygate4sd3_1
Xhold615 u_usb_cdc.u_sie.rx_valid VPWR VGND net934 sg13g2_dlygate4sd3_1
X_4493_ net702 VGND VPWR _0410_ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
X_3513_ _1455_ VPWR _0301_ VGND _1439_ _1456_ sg13g2_o21ai_1
X_3444_ net435 net581 _1408_ VPWR VGND sg13g2_nor2_1
Xhold637 _0313_ VPWR VGND net956 sg13g2_dlygate4sd3_1
Xhold648 u_usb_cdc.u_sie.crc16_q\[10\] VPWR VGND net967 sg13g2_dlygate4sd3_1
Xhold659 _0159_ VPWR VGND net978 sg13g2_dlygate4sd3_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_3375_ _1283_ net820 net814 _1364_ VPWR VGND sg13g2_a21o_1
X_2326_ _0558_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\] net809
+ VPWR VGND sg13g2_nand2b_1
X_2257_ _0487_ _0486_ _0489_ VPWR VGND sg13g2_xor2_1
XFILLER_27_28 VPWR VGND sg13g2_decap_8
X_2188_ u_usb_cdc.u_sie.u_phy_rx.rx_en_q _2040_ _2042_ VPWR VGND sg13g2_and2_1
XFILLER_4_128 VPWR VGND sg13g2_fill_1
XFILLER_0_323 VPWR VGND sg13g2_decap_8
XFILLER_49_828 VPWR VGND sg13g2_decap_8
XFILLER_17_703 VPWR VGND sg13g2_fill_1
XFILLER_1_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_32_706 VPWR VGND sg13g2_fill_2
XFILLER_8_412 VPWR VGND sg13g2_fill_1
XFILLER_40_772 VPWR VGND sg13g2_fill_2
XFILLER_12_485 VPWR VGND sg13g2_fill_2
XFILLER_9_957 VPWR VGND sg13g2_decap_4
XFILLER_4_662 VPWR VGND sg13g2_fill_1
XFILLER_4_651 VPWR VGND sg13g2_decap_8
X_3160_ _1205_ VPWR _0199_ VGND _1178_ _1204_ sg13g2_o21ai_1
X_2111_ _1968_ net890 VPWR VGND sg13g2_inv_2
X_3091_ _1152_ VPWR _0175_ VGND net828 _1160_ sg13g2_o21ai_1
Xhold1 u_usb_cdc.u_sie.u_phy_rx.dn_q\[2\] VPWR VGND net44 sg13g2_dlygate4sd3_1
XFILLER_48_850 VPWR VGND sg13g2_decap_8
X_3993_ net904 net709 _1828_ VPWR VGND sg13g2_nor2_1
XFILLER_22_238 VPWR VGND sg13g2_fill_2
X_2944_ net535 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ _1077_ _0111_ VPWR VGND sg13g2_mux2_1
X_2875_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net461 _1036_ _0083_ VPWR VGND sg13g2_mux2_1
Xhold401 _0087_ VPWR VGND net444 sg13g2_dlygate4sd3_1
Xhold445 u_usb_cdc.u_sie.data_q\[0\] VPWR VGND net488 sg13g2_dlygate4sd3_1
Xhold423 _0392_ VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold412 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[5\] VPWR VGND
+ net455 sg13g2_dlygate4sd3_1
Xhold434 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[63\] VPWR VGND
+ net477 sg13g2_dlygate4sd3_1
Xhold456 u_usb_cdc.u_ctrl_endp.addr_dd\[0\] VPWR VGND net499 sg13g2_dlygate4sd3_1
X_4476_ net729 VGND VPWR net188 u_usb_cdc.u_sie.rx_data\[0\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_1
Xhold478 _0112_ VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold467 _0114_ VPWR VGND net510 sg13g2_dlygate4sd3_1
Xhold489 u_usb_cdc.u_sie.u_phy_rx.dn_q\[0\] VPWR VGND net532 sg13g2_dlygate4sd3_1
X_3427_ net900 net435 _1397_ _0274_ VPWR VGND sg13g2_mux2_1
X_3358_ _1353_ net824 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[15\]
+ VPWR VGND sg13g2_nand2b_1
X_2309_ _0541_ net791 net788 VPWR VGND sg13g2_nand2_1
XFILLER_46_809 VPWR VGND sg13g2_decap_8
X_3289_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[24\] net821
+ _1291_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_599 VPWR VGND sg13g2_fill_2
XFILLER_16_1025 VPWR VGND sg13g2_decap_4
XFILLER_22_783 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_37_clk_regs clknet_3_5__leaf_clk_regs clknet_leaf_37_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_1_643 VPWR VGND sg13g2_decap_8
XFILLER_49_625 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_fill_2
XFILLER_48_146 VPWR VGND sg13g2_fill_1
XFILLER_17_555 VPWR VGND sg13g2_fill_1
XFILLER_45_897 VPWR VGND sg13g2_decap_8
XFILLER_32_558 VPWR VGND sg13g2_fill_2
XFILLER_13_750 VPWR VGND sg13g2_fill_1
X_2660_ _0869_ _0571_ _0868_ net596 net846 VPWR VGND sg13g2_a22oi_1
X_2591_ _0679_ net411 _0811_ _0000_ VPWR VGND sg13g2_a21o_1
X_4330_ net652 VGND VPWR net966 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[3\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_2
X_4261_ net657 VGND VPWR net335 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[23\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_3212_ _1233_ VPWR _0223_ VGND net723 net604 sg13g2_o21ai_1
X_4192_ net669 VGND VPWR net197 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[38\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_3143_ _1196_ VPWR _0191_ VGND net723 net605 sg13g2_o21ai_1
X_3074_ _1147_ VPWR _0171_ VGND _1915_ net634 sg13g2_o21ai_1
XFILLER_47_190 VPWR VGND sg13g2_fill_2
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_23_569 VPWR VGND sg13g2_decap_8
X_3976_ _1816_ VPWR _0404_ VGND _1951_ net613 sg13g2_o21ai_1
X_2927_ _1069_ net94 _1060_ VPWR VGND sg13g2_nand2_1
X_2858_ _1029_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[2\] _1028_
+ VPWR VGND sg13g2_xnor2_1
Xhold220 _0072_ VPWR VGND net263 sg13g2_dlygate4sd3_1
X_2789_ net638 _0955_ _0966_ VPWR VGND net771 sg13g2_nand3b_1
Xhold253 net20 VPWR VGND net296 sg13g2_dlygate4sd3_1
Xhold242 _1814_ VPWR VGND net285 sg13g2_dlygate4sd3_1
Xhold231 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[17\] VPWR VGND net274 sg13g2_dlygate4sd3_1
Xhold264 _0044_ VPWR VGND net307 sg13g2_dlygate4sd3_1
Xfanout700 net704 net700 VPWR VGND sg13g2_buf_8
Xhold275 _0215_ VPWR VGND net318 sg13g2_dlygate4sd3_1
XFILLER_49_26 VPWR VGND sg13g2_decap_8
Xhold286 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[4\] VPWR VGND net329 sg13g2_dlygate4sd3_1
X_4459_ net728 VGND VPWR net275 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[17\] clknet_leaf_25_clk_regs
+ sg13g2_dfrbpq_1
Xfanout722 _1911_ net722 VPWR VGND sg13g2_buf_8
Xfanout711 _1980_ net711 VPWR VGND sg13g2_buf_8
Xfanout733 net734 net733 VPWR VGND sg13g2_buf_8
Xhold297 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[10\] VPWR VGND net340 sg13g2_dlygate4sd3_1
Xfanout766 net560 net766 VPWR VGND sg13g2_buf_8
Xfanout755 net1043 net755 VPWR VGND sg13g2_buf_8
Xfanout744 net749 net744 VPWR VGND sg13g2_buf_8
Xfanout799 net800 net799 VPWR VGND sg13g2_buf_8
Xfanout788 net789 net788 VPWR VGND sg13g2_buf_8
Xfanout777 net778 net777 VPWR VGND sg13g2_buf_1
XFILLER_42_834 VPWR VGND sg13g2_fill_1
XFILLER_42_889 VPWR VGND sg13g2_decap_8
XFILLER_22_591 VPWR VGND sg13g2_fill_1
XFILLER_10_764 VPWR VGND sg13g2_fill_2
XFILLER_10_775 VPWR VGND sg13g2_fill_1
XFILLER_6_779 VPWR VGND sg13g2_fill_2
XFILLER_30_72 VPWR VGND sg13g2_fill_2
XFILLER_1_440 VPWR VGND sg13g2_decap_8
XFILLER_2_996 VPWR VGND sg13g2_decap_8
XFILLER_49_422 VPWR VGND sg13g2_decap_8
XFILLER_49_499 VPWR VGND sg13g2_decap_8
XFILLER_45_672 VPWR VGND sg13g2_fill_2
XFILLER_33_845 VPWR VGND sg13g2_fill_1
X_3830_ _0358_ _1713_ _1716_ _1703_ _1935_ VPWR VGND sg13g2_a22oi_1
X_3761_ _1661_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[70\] net628
+ VPWR VGND sg13g2_nand2_1
X_2712_ VGND VPWR _0911_ _0910_ _0909_ sg13g2_or2_1
X_3692_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[59\] net803 _1595_
+ VPWR VGND sg13g2_nor2b_1
X_2643_ _0847_ _0848_ _0846_ _0854_ VPWR VGND _0853_ sg13g2_nand4_1
X_2574_ _0676_ net622 _0662_ _0799_ VPWR VGND sg13g2_nand3_1
X_4313_ net652 VGND VPWR _0242_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\]
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
X_4244_ net656 VGND VPWR net256 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[6\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
XFILLER_19_18 VPWR VGND sg13g2_fill_2
XFILLER_28_606 VPWR VGND sg13g2_decap_8
X_4175_ net664 VGND VPWR net73 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[21\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
X_3126_ VGND VPWR net632 _1184_ _0186_ _1183_ sg13g2_a21oi_1
X_3057_ _1137_ net419 _1135_ VPWR VGND sg13g2_nand2_1
X_3959_ VGND VPWR net746 _0943_ _0395_ _1808_ sg13g2_a21oi_1
XFILLER_13_1017 VPWR VGND sg13g2_decap_8
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_738 VPWR VGND sg13g2_decap_4
XFILLER_47_915 VPWR VGND sg13g2_decap_8
Xfanout585 net587 net585 VPWR VGND sg13g2_buf_8
Xfanout596 net599 net596 VPWR VGND sg13g2_buf_8
XFILLER_26_160 VPWR VGND sg13g2_decap_4
XFILLER_42_631 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_52_clk_regs clknet_3_1__leaf_clk_regs clknet_leaf_52_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_41_163 VPWR VGND sg13g2_fill_2
XFILLER_44_7 VPWR VGND sg13g2_fill_2
X_2290_ net750 net752 net596 _0522_ VPWR VGND sg13g2_nor3_2
XFILLER_2_782 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_2_43 VPWR VGND sg13g2_fill_2
XFILLER_38_959 VPWR VGND sg13g2_decap_4
XFILLER_46_981 VPWR VGND sg13g2_decap_8
XFILLER_17_160 VPWR VGND sg13g2_fill_2
XFILLER_17_193 VPWR VGND sg13g2_fill_1
XFILLER_36_1028 VPWR VGND sg13g2_fill_1
X_3813_ net593 _0600_ _0512_ _1703_ VPWR VGND _1702_ sg13g2_nand4_1
XFILLER_33_675 VPWR VGND sg13g2_fill_2
X_3744_ net808 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[37\] _1645_
+ VPWR VGND sg13g2_nor2_1
X_3675_ VGND VPWR net802 _1578_ _1579_ _1923_ sg13g2_a21oi_1
X_2626_ net589 VPWR _0839_ VGND _0837_ _0838_ sg13g2_o21ai_1
X_2557_ _0783_ VPWR _0784_ VGND net622 _0766_ sg13g2_o21ai_1
X_2488_ net492 _0712_ _0715_ _0716_ VPWR VGND sg13g2_or3_1
X_4227_ net678 VGND VPWR net863 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[2\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
XFILLER_44_907 VPWR VGND sg13g2_decap_8
XFILLER_29_959 VPWR VGND sg13g2_decap_8
X_4158_ net663 VGND VPWR net444 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[4\]
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
X_3109_ _1171_ VPWR _0181_ VGND net827 _1172_ sg13g2_o21ai_1
X_4089_ net647 _1905_ net749 _1906_ VPWR VGND sg13g2_nand3_1
XFILLER_37_992 VPWR VGND sg13g2_decap_8
XFILLER_12_837 VPWR VGND sg13g2_fill_2
XFILLER_12_815 VPWR VGND sg13g2_fill_2
XFILLER_8_808 VPWR VGND sg13g2_fill_2
XFILLER_3_568 VPWR VGND sg13g2_fill_2
XFILLER_47_712 VPWR VGND sg13g2_decap_8
XFILLER_47_789 VPWR VGND sg13g2_decap_8
XFILLER_43_940 VPWR VGND sg13g2_decap_8
XFILLER_27_491 VPWR VGND sg13g2_fill_2
XFILLER_14_196 VPWR VGND sg13g2_fill_2
Xinput13 usb_dp_rx_i net13 VPWR VGND sg13g2_buf_1
XFILLER_6_340 VPWR VGND sg13g2_fill_1
XFILLER_6_384 VPWR VGND sg13g2_fill_1
X_3460_ _0661_ net622 _0751_ _1417_ VPWR VGND sg13g2_nor3_1
X_2411_ _0611_ _0616_ _0630_ _0641_ VGND VPWR _0640_ sg13g2_nor4_2
XFILLER_42_4 VPWR VGND sg13g2_fill_2
X_3391_ _1375_ VPWR _1376_ VGND net575 _1133_ sg13g2_o21ai_1
X_2342_ _0573_ VPWR _0574_ VGND net141 net601 sg13g2_o21ai_1
X_2273_ _0505_ _0486_ _0493_ VPWR VGND sg13g2_xnor2_1
X_4012_ _1843_ _1844_ _0518_ _1845_ VPWR VGND sg13g2_nand3_1
XFILLER_38_723 VPWR VGND sg13g2_fill_1
XFILLER_37_200 VPWR VGND sg13g2_fill_1
XFILLER_21_612 VPWR VGND sg13g2_fill_2
XFILLER_34_973 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
X_3727_ VGND VPWR _0647_ _0674_ _1629_ _0537_ sg13g2_a21oi_1
X_3658_ net602 VPWR _1563_ VGND net284 _1523_ sg13g2_o21ai_1
X_3589_ _1496_ _1968_ _1494_ VPWR VGND sg13g2_xnor2_1
X_2609_ _0619_ _0612_ _0827_ VPWR VGND _0613_ sg13g2_nand3b_1
XFILLER_0_505 VPWR VGND sg13g2_decap_8
XFILLER_28_255 VPWR VGND sg13g2_fill_1
XFILLER_28_277 VPWR VGND sg13g2_decap_8
XFILLER_40_921 VPWR VGND sg13g2_decap_4
XFILLER_40_943 VPWR VGND sg13g2_decap_8
XFILLER_11_188 VPWR VGND sg13g2_fill_2
Xheichips25_usb_cdc_36 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_3_365 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_26_1016 VPWR VGND sg13g2_decap_8
XFILLER_26_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_564 VPWR VGND sg13g2_fill_1
X_2960_ _1087_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2891_ _1038_ VPWR _0091_ VGND _1040_ net620 sg13g2_o21ai_1
XFILLER_42_280 VPWR VGND sg13g2_fill_1
Xhold616 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[1\] VPWR VGND
+ net935 sg13g2_dlygate4sd3_1
Xhold627 u_usb_cdc.u_ctrl_endp.in_dir_q VPWR VGND net946 sg13g2_dlygate4sd3_1
Xhold605 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[1\] VPWR VGND net924 sg13g2_dlygate4sd3_1
X_4492_ net733 VGND VPWR net12 u_usb_cdc.u_sie.u_phy_rx.dn_q\[2\] clknet_leaf_30_clk_regs
+ sg13g2_dfrbpq_1
X_3512_ _1456_ net562 _1453_ VPWR VGND sg13g2_xnor2_1
Xhold638 u_usb_cdc.u_ctrl_endp.req_q\[7\] VPWR VGND net957 sg13g2_dlygate4sd3_1
X_3443_ VGND VPWR _1914_ net581 _0280_ _1407_ sg13g2_a21oi_1
Xhold649 u_usb_cdc.u_ctrl_endp.state_q\[2\] VPWR VGND net968 sg13g2_dlygate4sd3_1
X_3374_ net814 _1283_ net820 _1363_ VPWR VGND sg13g2_nand3_1
X_2325_ _0557_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[3\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\] VPWR VGND sg13g2_nand2b_1
X_2256_ _0488_ _0486_ _0487_ VPWR VGND sg13g2_xnor2_1
X_2187_ _2041_ net53 net567 VPWR VGND sg13g2_nand2b_1
XFILLER_25_236 VPWR VGND sg13g2_decap_4
XFILLER_34_792 VPWR VGND sg13g2_fill_2
XFILLER_0_302 VPWR VGND sg13g2_decap_8
XFILLER_49_807 VPWR VGND sg13g2_decap_8
XFILLER_0_379 VPWR VGND sg13g2_decap_8
XFILLER_29_564 VPWR VGND sg13g2_fill_2
XFILLER_17_726 VPWR VGND sg13g2_fill_2
XFILLER_12_497 VPWR VGND sg13g2_decap_8
XFILLER_4_630 VPWR VGND sg13g2_fill_2
X_2110_ VPWR _1967_ net973 VGND sg13g2_inv_1
X_3090_ net832 _1159_ net764 _1160_ VPWR VGND sg13g2_nand3_1
Xhold2 u_usb_cdc.rstn_sq\[1\] VPWR VGND net45 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk_regs clknet_3_3__leaf_clk_regs clknet_leaf_7_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_16_770 VPWR VGND sg13g2_decap_8
X_3992_ VGND VPWR _1823_ _1826_ _1827_ _1822_ sg13g2_a21oi_1
XFILLER_35_567 VPWR VGND sg13g2_fill_2
XFILLER_35_589 VPWR VGND sg13g2_fill_2
XFILLER_16_781 VPWR VGND sg13g2_fill_1
X_2943_ net528 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ _1077_ _0110_ VPWR VGND sg13g2_mux2_1
X_2874_ _1036_ net740 _1035_ VPWR VGND sg13g2_nand2_2
Xhold402 net22 VPWR VGND net445 sg13g2_dlygate4sd3_1
Xhold424 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[59\] VPWR VGND
+ net467 sg13g2_dlygate4sd3_1
Xhold413 _0088_ VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold435 _0146_ VPWR VGND net478 sg13g2_dlygate4sd3_1
Xhold446 _0055_ VPWR VGND net489 sg13g2_dlygate4sd3_1
Xhold457 u_usb_cdc.u_ctrl_endp.endp_q\[3\] VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold468 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[25\] VPWR VGND
+ net511 sg13g2_dlygate4sd3_1
X_4475_ net732 VGND VPWR net451 u_usb_cdc.u_sie.u_phy_rx.rx_valid_q clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_1
Xhold479 u_usb_cdc.u_ctrl_endp.req_q\[11\] VPWR VGND net522 sg13g2_dlygate4sd3_1
X_3426_ net878 net473 _1397_ _0273_ VPWR VGND sg13g2_mux2_1
X_3357_ net824 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[39\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[47\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[55\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[63\] net817 _1352_
+ VPWR VGND sg13g2_mux4_1
X_2308_ net793 net789 _0540_ VPWR VGND sg13g2_and2_1
X_3288_ net823 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[16\]
+ _1290_ VPWR VGND sg13g2_nor2_1
X_2239_ _0471_ _0468_ _0470_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_718 VPWR VGND sg13g2_decap_8
XFILLER_26_567 VPWR VGND sg13g2_decap_8
XFILLER_22_740 VPWR VGND sg13g2_decap_4
XFILLER_5_416 VPWR VGND sg13g2_fill_2
XFILLER_1_622 VPWR VGND sg13g2_decap_8
XFILLER_49_604 VPWR VGND sg13g2_decap_8
XFILLER_1_699 VPWR VGND sg13g2_decap_8
XFILLER_45_876 VPWR VGND sg13g2_decap_8
XFILLER_44_342 VPWR VGND sg13g2_fill_1
XFILLER_32_548 VPWR VGND sg13g2_fill_1
X_2590_ _0048_ _0712_ _0758_ _0759_ _0811_ VPWR VGND sg13g2_nor4_1
X_4260_ net649 VGND VPWR net346 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[22\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
XFILLER_5_76 VPWR VGND sg13g2_fill_1
X_3211_ _1233_ net224 net604 VPWR VGND sg13g2_nand2_1
X_4191_ net668 VGND VPWR net114 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[37\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_3142_ _1196_ net172 net606 VPWR VGND sg13g2_nand2_1
X_3073_ _1147_ net304 net634 VPWR VGND sg13g2_nand2_1
XFILLER_36_887 VPWR VGND sg13g2_fill_1
X_3975_ _1816_ net266 net613 VPWR VGND sg13g2_nand2_1
X_2926_ _1067_ VPWR _0102_ VGND net618 _1068_ sg13g2_o21ai_1
X_2857_ _1028_ net1025 _1015_ VPWR VGND sg13g2_xnor2_1
X_2788_ _0965_ net742 _0964_ VPWR VGND sg13g2_nand2_1
Xhold210 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[50\] VPWR VGND
+ net253 sg13g2_dlygate4sd3_1
Xhold243 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[5\] VPWR VGND
+ net286 sg13g2_dlygate4sd3_1
Xhold221 net26 VPWR VGND net264 sg13g2_dlygate4sd3_1
Xhold232 _0387_ VPWR VGND net275 sg13g2_dlygate4sd3_1
Xhold254 _0244_ VPWR VGND net297 sg13g2_dlygate4sd3_1
Xhold265 _0058_ VPWR VGND net308 sg13g2_dlygate4sd3_1
X_4458_ net727 VGND VPWR _0386_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] clknet_leaf_25_clk_regs
+ sg13g2_dfrbpq_2
Xhold276 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[13\] VPWR VGND net319 sg13g2_dlygate4sd3_1
Xhold287 _0364_ VPWR VGND net330 sg13g2_dlygate4sd3_1
Xfanout723 _1910_ net723 VPWR VGND sg13g2_buf_8
X_3409_ net418 net578 _1391_ VPWR VGND sg13g2_nor2_1
Xfanout701 net704 net701 VPWR VGND sg13g2_buf_8
Xfanout712 _1980_ net712 VPWR VGND sg13g2_buf_1
Xhold298 _0380_ VPWR VGND net341 sg13g2_dlygate4sd3_1
Xfanout734 net737 net734 VPWR VGND sg13g2_buf_8
Xfanout767 net488 net767 VPWR VGND sg13g2_buf_8
Xfanout756 net1043 net756 VPWR VGND sg13g2_buf_2
Xfanout745 net746 net745 VPWR VGND sg13g2_buf_8
X_4389_ net698 VGND VPWR net432 u_usb_cdc.u_sie.delay_cnt_q\[1\] clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_2
Xfanout789 net790 net789 VPWR VGND sg13g2_buf_1
Xfanout778 net1021 net778 VPWR VGND sg13g2_buf_8
XFILLER_39_681 VPWR VGND sg13g2_decap_8
XFILLER_14_537 VPWR VGND sg13g2_decap_4
XFILLER_14_63 VPWR VGND sg13g2_fill_2
XFILLER_2_920 VPWR VGND sg13g2_fill_2
XFILLER_1_430 VPWR VGND sg13g2_decap_4
XFILLER_2_975 VPWR VGND sg13g2_decap_8
XFILLER_49_401 VPWR VGND sg13g2_decap_8
XFILLER_49_478 VPWR VGND sg13g2_decap_8
XFILLER_45_684 VPWR VGND sg13g2_decap_8
X_3760_ _1637_ VPWR _0344_ VGND _1659_ _1660_ sg13g2_o21ai_1
X_2711_ VGND VPWR _0910_ _2047_ _1975_ sg13g2_or2_1
X_3691_ net799 _1592_ _1593_ _1594_ VPWR VGND sg13g2_nor3_1
X_2642_ _0849_ _0850_ _0851_ _0852_ _0853_ VPWR VGND sg13g2_nor4_1
X_2573_ _0798_ _0673_ _0769_ VPWR VGND sg13g2_nand2_1
X_4312_ net657 VGND VPWR _0241_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[2\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_2
X_4243_ net673 VGND VPWR net287 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[5\]
+ clknet_leaf_47_clk_regs sg13g2_dfrbpq_1
X_4174_ net662 VGND VPWR net95 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[20\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
X_3125_ _1184_ net760 _1141_ VPWR VGND sg13g2_nand2_1
X_3056_ VGND VPWR _1986_ _1135_ _0164_ _1136_ sg13g2_a21oi_1
X_3958_ net751 net746 _1808_ VPWR VGND sg13g2_nor2_1
X_2909_ _1055_ VPWR _0097_ VGND net619 _1056_ sg13g2_o21ai_1
X_3889_ _1758_ VPWR _0374_ VGND net348 _1759_ sg13g2_o21ai_1
XFILLER_3_717 VPWR VGND sg13g2_decap_8
XFILLER_2_205 VPWR VGND sg13g2_fill_2
XFILLER_2_238 VPWR VGND sg13g2_fill_1
Xfanout586 net587 net586 VPWR VGND sg13g2_buf_1
Xfanout597 net599 net597 VPWR VGND sg13g2_buf_8
XFILLER_18_128 VPWR VGND sg13g2_fill_1
XFILLER_15_879 VPWR VGND sg13g2_decap_8
XFILLER_30_838 VPWR VGND sg13g2_fill_2
XFILLER_41_153 VPWR VGND sg13g2_fill_1
XFILLER_10_584 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_21_clk_regs clknet_3_6__leaf_clk_regs clknet_leaf_21_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_6_555 VPWR VGND sg13g2_fill_1
XFILLER_1_260 VPWR VGND sg13g2_fill_1
XFILLER_37_7 VPWR VGND sg13g2_decap_4
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_2_99 VPWR VGND sg13g2_fill_1
XFILLER_46_960 VPWR VGND sg13g2_decap_8
XFILLER_36_1007 VPWR VGND sg13g2_decap_8
X_3812_ _1702_ _1701_ _1972_ _2017_ net848 VPWR VGND sg13g2_a22oi_1
X_3743_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[45\] net805 _1644_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_9_393 VPWR VGND sg13g2_decap_8
X_3674_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[50\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[58\]
+ net807 _1578_ VPWR VGND sg13g2_mux2_1
X_2625_ _1928_ _0624_ _0838_ VPWR VGND sg13g2_nor2_1
X_2556_ _0774_ _0776_ _0780_ _0782_ _0783_ VPWR VGND sg13g2_nor4_1
X_2487_ _0715_ net641 _0714_ VPWR VGND sg13g2_nand2_1
X_4226_ net681 VGND VPWR net860 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[1\]
+ clknet_leaf_20_clk_regs sg13g2_dfrbpq_1
X_4157_ net661 VGND VPWR net434 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[3\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
XFILLER_29_938 VPWR VGND sg13g2_decap_8
X_3108_ net830 _1159_ net758 _1172_ VPWR VGND sg13g2_nand3_1
X_4088_ _1905_ net547 _1031_ VPWR VGND sg13g2_nand2_1
X_3039_ _1025_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[1\] _1031_
+ _1129_ VPWR VGND sg13g2_mux2_1
XFILLER_23_153 VPWR VGND sg13g2_decap_4
XFILLER_3_547 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1016 VPWR VGND sg13g2_decap_8
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_234 VPWR VGND sg13g2_fill_2
XFILLER_47_768 VPWR VGND sg13g2_decap_8
XFILLER_15_621 VPWR VGND sg13g2_fill_1
XFILLER_28_993 VPWR VGND sg13g2_decap_8
XFILLER_46_278 VPWR VGND sg13g2_fill_1
XFILLER_43_996 VPWR VGND sg13g2_decap_8
XFILLER_15_665 VPWR VGND sg13g2_decap_4
XFILLER_30_635 VPWR VGND sg13g2_decap_8
XFILLER_11_860 VPWR VGND sg13g2_decap_8
XFILLER_10_392 VPWR VGND sg13g2_decap_4
X_2410_ _0640_ net743 _0638_ VPWR VGND sg13g2_nand2_2
X_3390_ _1375_ _1133_ _1374_ VPWR VGND sg13g2_nand2_1
X_2341_ _0573_ _0568_ _0571_ VPWR VGND sg13g2_nand2_1
X_2272_ u_usb_cdc.u_sie.crc16_q\[5\] u_usb_cdc.u_sie.crc16_q\[4\] u_usb_cdc.u_sie.crc16_q\[7\]
+ u_usb_cdc.u_sie.crc16_q\[6\] _0504_ VPWR VGND sg13g2_nor4_1
XFILLER_42_1022 VPWR VGND sg13g2_decap_8
X_4011_ _1844_ _1966_ net837 net765 net842 VPWR VGND sg13g2_a22oi_1
XFILLER_37_212 VPWR VGND sg13g2_fill_1
XFILLER_20_112 VPWR VGND sg13g2_fill_2
X_3726_ net773 VPWR _1628_ VGND _0543_ _0657_ sg13g2_o21ai_1
X_3657_ VPWR VGND net637 net627 _1561_ _1499_ _1562_ _1552_ sg13g2_a221oi_1
X_3588_ _0337_ net579 _1969_ net583 _1954_ VPWR VGND sg13g2_a22oi_1
X_2608_ _0826_ VPWR _0011_ VGND _1927_ _0817_ sg13g2_o21ai_1
X_2539_ VGND VPWR _0671_ _0765_ _0766_ _0764_ sg13g2_a21oi_1
X_4209_ net670 VGND VPWR net151 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[55\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
XFILLER_17_908 VPWR VGND sg13g2_fill_2
XFILLER_44_727 VPWR VGND sg13g2_fill_1
XFILLER_44_716 VPWR VGND sg13g2_fill_1
XFILLER_24_484 VPWR VGND sg13g2_decap_8
XFILLER_8_617 VPWR VGND sg13g2_fill_2
XFILLER_8_628 VPWR VGND sg13g2_fill_1
XFILLER_40_999 VPWR VGND sg13g2_decap_8
XFILLER_8_639 VPWR VGND sg13g2_fill_2
Xheichips25_usb_cdc_37 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_16_930 VPWR VGND sg13g2_decap_4
XFILLER_15_484 VPWR VGND sg13g2_decap_8
XFILLER_42_270 VPWR VGND sg13g2_fill_1
X_2890_ VGND VPWR _1044_ _1042_ _1041_ sg13g2_or2_1
XFILLER_31_988 VPWR VGND sg13g2_decap_8
Xhold617 _0252_ VPWR VGND net936 sg13g2_dlygate4sd3_1
Xhold606 _0928_ VPWR VGND net925 sg13g2_dlygate4sd3_1
X_4491_ net733 VGND VPWR net44 u_usb_cdc.u_sie.u_phy_rx.dn_q\[1\] clknet_leaf_30_clk_regs
+ sg13g2_dfrbpq_1
X_3511_ _1455_ net562 _1437_ VPWR VGND sg13g2_nand2_1
Xhold639 _0008_ VPWR VGND net958 sg13g2_dlygate4sd3_1
X_3442_ net473 net581 _1407_ VPWR VGND sg13g2_nor2_1
Xhold628 _0836_ VPWR VGND net947 sg13g2_dlygate4sd3_1
X_3373_ net629 _1362_ _0255_ VPWR VGND sg13g2_nor2_1
X_2324_ VGND VPWR _0555_ _0556_ _0554_ _0549_ sg13g2_a21oi_2
X_2255_ u_usb_cdc.u_sie.data_q\[3\] net913 _0487_ VPWR VGND sg13g2_xor2_1
X_2186_ net567 net53 _2040_ VPWR VGND sg13g2_nor2b_2
XFILLER_26_705 VPWR VGND sg13g2_fill_2
XFILLER_38_576 VPWR VGND sg13g2_fill_2
XFILLER_38_598 VPWR VGND sg13g2_decap_4
XFILLER_33_281 VPWR VGND sg13g2_decap_4
X_3709_ _1612_ net1005 net597 VPWR VGND sg13g2_nand2_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_1017 VPWR VGND sg13g2_decap_8
XFILLER_1_804 VPWR VGND sg13g2_decap_8
XFILLER_0_358 VPWR VGND sg13g2_decap_8
XFILLER_44_513 VPWR VGND sg13g2_decap_4
XFILLER_16_226 VPWR VGND sg13g2_fill_2
XFILLER_17_52 VPWR VGND sg13g2_fill_1
XFILLER_32_708 VPWR VGND sg13g2_fill_1
XFILLER_9_926 VPWR VGND sg13g2_fill_1
XFILLER_13_977 VPWR VGND sg13g2_fill_1
XFILLER_12_487 VPWR VGND sg13g2_fill_1
XFILLER_32_1010 VPWR VGND sg13g2_decap_8
XFILLER_0_881 VPWR VGND sg13g2_decap_8
Xhold3 u_usb_cdc.u_sie.u_phy_rx.dp_q\[2\] VPWR VGND net46 sg13g2_dlygate4sd3_1
XFILLER_48_885 VPWR VGND sg13g2_decap_8
X_3991_ _1824_ _1825_ _1705_ _1826_ VPWR VGND sg13g2_nand3_1
X_2942_ net537 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ _1077_ _0109_ VPWR VGND sg13g2_mux2_1
X_2873_ _1985_ _1019_ _1035_ VPWR VGND sg13g2_and2_1
XFILLER_8_992 VPWR VGND sg13g2_decap_8
Xhold403 _1313_ VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold425 _0142_ VPWR VGND net468 sg13g2_dlygate4sd3_1
Xhold436 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[62\] VPWR VGND
+ net479 sg13g2_dlygate4sd3_1
Xhold414 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[8\] VPWR VGND net457 sg13g2_dlygate4sd3_1
Xhold469 _0108_ VPWR VGND net512 sg13g2_dlygate4sd3_1
Xhold447 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[2\] VPWR VGND
+ net490 sg13g2_dlygate4sd3_1
X_4474_ net689 VGND VPWR _0400_ u_usb_cdc.sie_in_data_ack clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_2
Xhold458 u_usb_cdc.u_sie.u_phy_rx.rx_eop_q VPWR VGND net501 sg13g2_dlygate4sd3_1
X_3425_ net897 net566 _1397_ _0272_ VPWR VGND sg13g2_mux2_1
X_3356_ _0249_ _1350_ _1351_ net616 _2012_ VPWR VGND sg13g2_a22oi_1
X_3287_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[0\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[8\]
+ net824 _1289_ VPWR VGND sg13g2_mux2_1
X_2307_ _0539_ net791 VPWR VGND net784 sg13g2_nand2b_2
X_2238_ _0470_ _0456_ _0469_ VPWR VGND sg13g2_xnor2_1
X_2169_ _2025_ net626 net625 VPWR VGND sg13g2_nand2_1
XFILLER_1_678 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_46_clk_regs clknet_3_4__leaf_clk_regs clknet_leaf_46_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_48_115 VPWR VGND sg13g2_decap_4
XFILLER_17_502 VPWR VGND sg13g2_fill_2
XFILLER_45_855 VPWR VGND sg13g2_decap_8
XFILLER_44_398 VPWR VGND sg13g2_fill_1
XFILLER_9_756 VPWR VGND sg13g2_fill_1
XFILLER_5_984 VPWR VGND sg13g2_decap_8
X_3210_ _1232_ net828 _1194_ VPWR VGND sg13g2_nand2_2
X_4190_ net668 VGND VPWR net206 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[36\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
X_3141_ _1195_ net711 _1194_ VPWR VGND sg13g2_nand2_1
X_3072_ _1146_ VPWR _0170_ VGND net720 net635 sg13g2_o21ai_1
XFILLER_36_844 VPWR VGND sg13g2_fill_2
XFILLER_48_682 VPWR VGND sg13g2_decap_8
XFILLER_39_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_1016 VPWR VGND sg13g2_decap_8
XFILLER_36_866 VPWR VGND sg13g2_fill_2
XFILLER_36_877 VPWR VGND sg13g2_fill_1
XFILLER_47_192 VPWR VGND sg13g2_fill_1
X_3974_ _1815_ VPWR _0403_ VGND _1948_ net613 sg13g2_o21ai_1
X_2925_ _1068_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net644 VPWR VGND sg13g2_nand2_1
X_2856_ VGND VPWR _1986_ _1025_ _1027_ _1017_ sg13g2_a21oi_1
X_2787_ _0963_ _0961_ _0964_ VPWR VGND sg13g2_nor2b_2
Xhold211 _0133_ VPWR VGND net254 sg13g2_dlygate4sd3_1
Xhold200 _0137_ VPWR VGND net243 sg13g2_dlygate4sd3_1
Xhold244 _0172_ VPWR VGND net287 sg13g2_dlygate4sd3_1
Xhold233 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[58\] VPWR
+ VGND net276 sg13g2_dlygate4sd3_1
Xhold222 _0250_ VPWR VGND net265 sg13g2_dlygate4sd3_1
XFILLER_46_1009 VPWR VGND sg13g2_decap_8
Xhold255 u_usb_cdc.sie_out_data\[4\] VPWR VGND net298 sg13g2_dlygate4sd3_1
Xhold266 _0418_ VPWR VGND net309 sg13g2_dlygate4sd3_1
Xhold277 _0383_ VPWR VGND net320 sg13g2_dlygate4sd3_1
X_4457_ net727 VGND VPWR _0385_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[15\] clknet_leaf_25_clk_regs
+ sg13g2_dfrbpq_1
Xfanout724 _1910_ net724 VPWR VGND sg13g2_buf_1
Xhold299 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[49\] VPWR
+ VGND net342 sg13g2_dlygate4sd3_1
Xhold288 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[19\] VPWR
+ VGND net331 sg13g2_dlygate4sd3_1
X_3408_ _1387_ _1389_ _1390_ VPWR VGND sg13g2_nor2_2
Xfanout702 net703 net702 VPWR VGND sg13g2_buf_8
Xfanout713 net715 net713 VPWR VGND sg13g2_buf_8
Xfanout735 net737 net735 VPWR VGND sg13g2_buf_8
Xfanout757 net1012 net757 VPWR VGND sg13g2_buf_8
X_4388_ net697 VGND VPWR net355 u_usb_cdc.u_sie.delay_cnt_q\[0\] clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_2
Xfanout746 net747 net746 VPWR VGND sg13g2_buf_1
X_3339_ VGND VPWR net822 _1999_ _1336_ _1286_ sg13g2_a21oi_1
Xfanout768 net769 net768 VPWR VGND sg13g2_buf_8
Xfanout779 net783 net779 VPWR VGND sg13g2_buf_8
XFILLER_46_619 VPWR VGND sg13g2_fill_2
XFILLER_14_505 VPWR VGND sg13g2_decap_8
XFILLER_10_766 VPWR VGND sg13g2_fill_1
XFILLER_5_236 VPWR VGND sg13g2_fill_2
XFILLER_30_41 VPWR VGND sg13g2_decap_4
XFILLER_2_954 VPWR VGND sg13g2_decap_8
XFILLER_7_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_49_457 VPWR VGND sg13g2_decap_8
XFILLER_18_811 VPWR VGND sg13g2_fill_1
XFILLER_45_674 VPWR VGND sg13g2_fill_1
XFILLER_13_571 VPWR VGND sg13g2_fill_1
X_2710_ _0909_ _2042_ _2035_ VPWR VGND sg13g2_nand2b_1
X_3690_ net803 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[35\] _1593_
+ VPWR VGND sg13g2_nor2_1
X_2641_ u_usb_cdc.u_sie.addr_q\[2\] u_usb_cdc.addr\[2\] _0852_ VPWR VGND sg13g2_xor2_1
X_2572_ u_usb_cdc.u_ctrl_endp.rec_q\[1\] _0641_ _1936_ _0797_ VPWR VGND net623 sg13g2_nand4_1
XFILLER_5_770 VPWR VGND sg13g2_fill_1
X_4311_ net652 VGND VPWR net893 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\]
+ clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
X_4242_ net672 VGND VPWR _0171_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[4\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_4173_ net665 VGND VPWR net249 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[19\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
X_3124_ net331 net632 _1183_ VPWR VGND sg13g2_nor2_1
X_3055_ net801 _1135_ _1136_ VPWR VGND sg13g2_nor2_1
XFILLER_24_803 VPWR VGND sg13g2_fill_1
XFILLER_11_519 VPWR VGND sg13g2_fill_2
X_3957_ net708 net976 _1807_ _0394_ VPWR VGND sg13g2_a21o_1
Xclkbuf_0_clk_regs clk_regs clknet_0_clk_regs VPWR VGND sg13g2_buf_8
X_2908_ _1056_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net645 VPWR VGND sg13g2_nand2_1
X_3888_ _1759_ net615 _1754_ VPWR VGND sg13g2_nand2_1
X_2839_ VPWR VGND u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\]
+ _2028_ _1909_ _1011_ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] sg13g2_a221oi_1
X_4509_ net729 VGND VPWR _0039_ u_usb_cdc.clk_cnt_q\[0\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
XFILLER_4_8 VPWR VGND sg13g2_decap_8
Xfanout587 _1002_ net587 VPWR VGND sg13g2_buf_8
Xfanout576 _1419_ net576 VPWR VGND sg13g2_buf_2
Xfanout598 net599 net598 VPWR VGND sg13g2_buf_1
XFILLER_27_630 VPWR VGND sg13g2_fill_1
XFILLER_27_674 VPWR VGND sg13g2_fill_1
XFILLER_26_184 VPWR VGND sg13g2_fill_1
XFILLER_41_165 VPWR VGND sg13g2_fill_1
XFILLER_6_512 VPWR VGND sg13g2_decap_8
XFILLER_6_578 VPWR VGND sg13g2_decap_8
XFILLER_6_589 VPWR VGND sg13g2_fill_2
XFILLER_29_1015 VPWR VGND sg13g2_decap_8
XFILLER_2_740 VPWR VGND sg13g2_decap_4
XFILLER_44_9 VPWR VGND sg13g2_fill_1
XFILLER_2_67 VPWR VGND sg13g2_fill_2
XFILLER_2_78 VPWR VGND sg13g2_fill_1
XFILLER_33_644 VPWR VGND sg13g2_fill_2
X_3811_ net841 net847 _1701_ VPWR VGND sg13g2_nor2_2
XFILLER_33_677 VPWR VGND sg13g2_fill_1
XFILLER_21_828 VPWR VGND sg13g2_fill_2
X_3742_ _1642_ VPWR _1643_ VGND net798 _1640_ sg13g2_o21ai_1
X_3673_ _1576_ VPWR _1577_ VGND net807 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[34\]
+ sg13g2_o21ai_1
X_2624_ _1918_ _1929_ _0549_ _0837_ VPWR VGND sg13g2_nor3_1
X_2555_ _0781_ VPWR _0782_ VGND _0684_ _0686_ sg13g2_o21ai_1
X_2486_ net756 _0602_ _0714_ VPWR VGND sg13g2_nor2_2
X_4225_ net678 VGND VPWR net138 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[71\]
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
X_4156_ net661 VGND VPWR net491 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[2\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_1
XFILLER_29_917 VPWR VGND sg13g2_decap_8
X_3107_ _1171_ net222 _1151_ VPWR VGND sg13g2_nand2_1
X_4087_ net884 _1904_ _1128_ _0427_ VPWR VGND sg13g2_mux2_1
X_3038_ VGND VPWR _1127_ _1128_ _0593_ _0592_ sg13g2_a21oi_2
XFILLER_24_655 VPWR VGND sg13g2_decap_4
XFILLER_12_817 VPWR VGND sg13g2_fill_1
XFILLER_24_666 VPWR VGND sg13g2_fill_2
XFILLER_12_839 VPWR VGND sg13g2_fill_1
XFILLER_11_349 VPWR VGND sg13g2_fill_1
XFILLER_47_747 VPWR VGND sg13g2_decap_8
XFILLER_46_246 VPWR VGND sg13g2_decap_4
XFILLER_28_972 VPWR VGND sg13g2_decap_8
XFILLER_42_430 VPWR VGND sg13g2_fill_1
XFILLER_43_975 VPWR VGND sg13g2_decap_8
XFILLER_14_198 VPWR VGND sg13g2_fill_1
XFILLER_42_496 VPWR VGND sg13g2_decap_4
XFILLER_7_865 VPWR VGND sg13g2_decap_4
X_2340_ _0572_ net594 _0570_ VPWR VGND sg13g2_nand2_1
XFILLER_42_1001 VPWR VGND sg13g2_decap_8
X_2271_ u_usb_cdc.u_sie.crc16_q\[3\] u_usb_cdc.u_sie.crc16_q\[2\] _0503_ VPWR VGND
+ sg13g2_nor2_1
X_4010_ _1843_ _1955_ net845 u_usb_cdc.u_sie.pid_q\[2\] net836 VPWR VGND sg13g2_a22oi_1
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_21_614 VPWR VGND sg13g2_fill_1
X_3725_ VGND VPWR _0545_ _0821_ _1627_ _1513_ sg13g2_a21oi_1
X_3656_ _1553_ VPWR _1561_ VGND net795 _1560_ sg13g2_o21ai_1
X_3587_ _0336_ net580 _1966_ net584 _1955_ VPWR VGND sg13g2_a22oi_1
X_2607_ _0617_ _0820_ net742 _0826_ VPWR VGND _0824_ sg13g2_nand4_1
X_2538_ u_usb_cdc.u_ctrl_endp.req_q\[4\] net851 u_usb_cdc.u_ctrl_endp.req_q\[7\] _0765_
+ VPWR VGND sg13g2_or3_1
X_2469_ net763 _0693_ _0697_ VPWR VGND sg13g2_nor2_1
X_4208_ net670 VGND VPWR net243 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[54\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_4139_ net687 VGND VPWR net263 u_usb_cdc.u_sie.addr_q\[0\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_19_1025 VPWR VGND sg13g2_decap_4
XFILLER_25_997 VPWR VGND sg13g2_decap_8
XFILLER_40_978 VPWR VGND sg13g2_decap_8
XFILLER_4_824 VPWR VGND sg13g2_fill_1
XFILLER_31_967 VPWR VGND sg13g2_decap_8
X_3510_ _1451_ VPWR _0300_ VGND _1439_ _1454_ sg13g2_o21ai_1
XFILLER_7_684 VPWR VGND sg13g2_decap_4
Xhold607 u_usb_cdc.u_ctrl_endp.max_length_q\[1\] VPWR VGND net926 sg13g2_dlygate4sd3_1
Xhold618 _0059_ VPWR VGND net937 sg13g2_dlygate4sd3_1
X_4490_ net733 VGND VPWR net48 u_usb_cdc.u_sie.u_phy_rx.dn_q\[0\] clknet_leaf_30_clk_regs
+ sg13g2_dfrbpq_1
X_3441_ VGND VPWR _1915_ net581 _0279_ _1406_ sg13g2_a21oi_1
Xhold629 _0016_ VPWR VGND net948 sg13g2_dlygate4sd3_1
X_3372_ _1362_ net820 _1283_ VPWR VGND sg13g2_xnor2_1
X_2323_ VGND VPWR _0555_ u_usb_cdc.u_ctrl_endp.state_q\[3\] net769 sg13g2_or2_1
X_2254_ _0486_ net920 u_usb_cdc.u_sie.data_q\[4\] VPWR VGND sg13g2_xnor2_1
XFILLER_38_500 VPWR VGND sg13g2_fill_1
X_2185_ _2037_ _2038_ _2035_ _2039_ VPWR VGND sg13g2_nand3_1
XFILLER_22_934 VPWR VGND sg13g2_fill_1
XFILLER_34_794 VPWR VGND sg13g2_fill_1
XFILLER_21_488 VPWR VGND sg13g2_fill_2
X_3708_ net602 VPWR _1611_ VGND net266 _1523_ sg13g2_o21ai_1
X_3639_ _0652_ VPWR _1544_ VGND net792 _0533_ sg13g2_o21ai_1
XFILLER_0_337 VPWR VGND sg13g2_decap_8
XFILLER_17_728 VPWR VGND sg13g2_fill_1
XFILLER_17_64 VPWR VGND sg13g2_decap_8
XFILLER_17_75 VPWR VGND sg13g2_fill_1
XFILLER_13_912 VPWR VGND sg13g2_fill_2
XFILLER_13_945 VPWR VGND sg13g2_fill_1
XFILLER_9_949 VPWR VGND sg13g2_decap_4
XFILLER_4_687 VPWR VGND sg13g2_fill_1
Xhold4 u_usb_cdc.u_sie.u_phy_rx.dp_q\[1\] VPWR VGND net47 sg13g2_dlygate4sd3_1
XFILLER_48_864 VPWR VGND sg13g2_decap_8
X_3990_ _1825_ _1968_ net837 _1953_ net845 VPWR VGND sg13g2_a22oi_1
X_2941_ net511 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ _1077_ _0108_ VPWR VGND sg13g2_mux2_1
XFILLER_30_252 VPWR VGND sg13g2_fill_2
XFILLER_30_263 VPWR VGND sg13g2_fill_1
X_2872_ net833 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ _1034_ VPWR VGND sg13g2_nor3_1
XFILLER_8_971 VPWR VGND sg13g2_decap_8
X_4473_ net736 VGND VPWR net534 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_2
Xhold404 _0246_ VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold426 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[58\] VPWR VGND
+ net469 sg13g2_dlygate4sd3_1
Xhold415 _0378_ VPWR VGND net458 sg13g2_dlygate4sd3_1
X_3424_ net923 net559 _1397_ _0271_ VPWR VGND sg13g2_mux2_1
Xhold448 _0085_ VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold459 _0945_ VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold437 _0145_ VPWR VGND net480 sg13g2_dlygate4sd3_1
X_3355_ VGND VPWR net166 net629 _1351_ net617 sg13g2_a21oi_1
X_3286_ VGND VPWR _1288_ net813 net814 sg13g2_or2_1
X_2306_ net772 _1926_ _0537_ _0538_ VPWR VGND sg13g2_nor3_1
X_2237_ _0469_ net763 net765 VPWR VGND sg13g2_xnor2_1
XFILLER_39_864 VPWR VGND sg13g2_fill_1
X_2168_ _2024_ net747 _2021_ VPWR VGND sg13g2_nand2_1
X_2099_ VPWR _1956_ net913 VGND sg13g2_inv_1
XFILLER_1_657 VPWR VGND sg13g2_decap_8
XFILLER_49_639 VPWR VGND sg13g2_decap_8
XFILLER_45_812 VPWR VGND sg13g2_fill_2
XFILLER_45_801 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk_regs clknet_3_2__leaf_clk_regs clknet_leaf_15_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_13_720 VPWR VGND sg13g2_decap_4
XFILLER_44_40 VPWR VGND sg13g2_fill_1
XFILLER_44_388 VPWR VGND sg13g2_fill_2
XFILLER_13_764 VPWR VGND sg13g2_fill_2
XFILLER_13_786 VPWR VGND sg13g2_fill_1
XFILLER_8_223 VPWR VGND sg13g2_fill_2
XFILLER_9_746 VPWR VGND sg13g2_decap_4
XFILLER_9_779 VPWR VGND sg13g2_fill_2
XFILLER_5_963 VPWR VGND sg13g2_decap_8
X_3140_ _1158_ _1193_ _1194_ VPWR VGND sg13g2_nor2_1
X_3071_ _1146_ net184 net635 VPWR VGND sg13g2_nand2_1
XFILLER_48_661 VPWR VGND sg13g2_decap_8
X_3973_ _1815_ net232 net613 VPWR VGND sg13g2_nand2_1
X_2924_ _1067_ net248 _1060_ VPWR VGND sg13g2_nand2_1
XFILLER_31_583 VPWR VGND sg13g2_decap_8
X_2855_ _1026_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[1\] _1025_
+ VPWR VGND sg13g2_nand2b_1
Xhold201 net24 VPWR VGND net244 sg13g2_dlygate4sd3_1
X_2786_ VGND VPWR _1971_ _0962_ _0963_ net851 sg13g2_a21oi_1
Xhold234 _0225_ VPWR VGND net277 sg13g2_dlygate4sd3_1
Xhold212 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[6\] VPWR VGND
+ net255 sg13g2_dlygate4sd3_1
Xhold223 u_usb_cdc.u_sie.rx_data\[3\] VPWR VGND net266 sg13g2_dlygate4sd3_1
Xhold245 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[2\] VPWR VGND
+ net288 sg13g2_dlygate4sd3_1
Xhold278 u_usb_cdc.u_sie.in_byte_q\[2\] VPWR VGND net321 sg13g2_dlygate4sd3_1
Xhold256 _0054_ VPWR VGND net299 sg13g2_dlygate4sd3_1
X_4456_ net727 VGND VPWR _0384_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[14\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
Xhold267 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[5\] VPWR VGND net310 sg13g2_dlygate4sd3_1
Xhold289 _0186_ VPWR VGND net332 sg13g2_dlygate4sd3_1
X_3407_ _1389_ net743 _1388_ VPWR VGND sg13g2_nand2_2
X_4387_ net699 VGND VPWR _0315_ u_usb_cdc.sie_in_req clknet_leaf_36_clk_regs sg13g2_dfrbpq_2
Xfanout703 net704 net703 VPWR VGND sg13g2_buf_8
Xfanout714 net715 net714 VPWR VGND sg13g2_buf_1
Xfanout736 net737 net736 VPWR VGND sg13g2_buf_2
Xfanout758 net1024 net758 VPWR VGND sg13g2_buf_8
X_3338_ VGND VPWR _1335_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[21\]
+ net823 sg13g2_or2_1
Xfanout747 net748 net747 VPWR VGND sg13g2_buf_8
Xfanout725 net738 net725 VPWR VGND sg13g2_buf_8
Xfanout769 u_usb_cdc.endp\[0\] net769 VPWR VGND sg13g2_buf_8
X_3269_ _1273_ net770 net940 VPWR VGND sg13g2_nand2_1
XFILLER_39_661 VPWR VGND sg13g2_decap_4
XFILLER_38_193 VPWR VGND sg13g2_fill_2
XFILLER_14_528 VPWR VGND sg13g2_decap_4
XFILLER_14_517 VPWR VGND sg13g2_fill_2
XFILLER_22_561 VPWR VGND sg13g2_fill_1
XFILLER_14_65 VPWR VGND sg13g2_fill_1
XFILLER_1_454 VPWR VGND sg13g2_decap_8
XFILLER_49_436 VPWR VGND sg13g2_decap_8
XFILLER_45_664 VPWR VGND sg13g2_decap_4
X_2640_ u_usb_cdc.u_sie.addr_q\[1\] u_usb_cdc.addr\[1\] _0851_ VPWR VGND sg13g2_xor2_1
XFILLER_9_598 VPWR VGND sg13g2_decap_8
X_2571_ VGND VPWR _0635_ _0662_ _0796_ _0620_ sg13g2_a21oi_1
XFILLER_5_782 VPWR VGND sg13g2_decap_8
X_4310_ net657 VGND VPWR _0239_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[0\]
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
X_4241_ net656 VGND VPWR _0170_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[3\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_4172_ net660 VGND VPWR net183 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[18\]
+ clknet_leaf_10_clk_regs sg13g2_dfrbpq_1
X_3123_ VGND VPWR net632 _1182_ _0185_ _1181_ sg13g2_a21oi_1
XFILLER_27_108 VPWR VGND sg13g2_fill_1
X_3054_ net809 net931 _1135_ _0163_ VPWR VGND sg13g2_mux2_1
XFILLER_36_653 VPWR VGND sg13g2_decap_8
X_3956_ _1978_ net368 net708 _1806_ _1807_ VPWR VGND sg13g2_nor4_1
X_2907_ _1055_ net220 _1037_ VPWR VGND sg13g2_nand2_1
X_3887_ _1758_ net348 _1755_ VPWR VGND sg13g2_nand2_1
X_2838_ _1010_ _1008_ net626 VPWR VGND sg13g2_nand2b_1
X_2769_ _0946_ _0479_ _0441_ _0947_ VPWR VGND sg13g2_a21o_1
X_4508_ net729 VGND VPWR _0041_ u_usb_cdc.clk_gate_q clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
X_4439_ net730 VGND VPWR net497 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[6\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_47_929 VPWR VGND sg13g2_decap_8
Xfanout577 _1419_ net577 VPWR VGND sg13g2_buf_1
Xfanout588 _0622_ net588 VPWR VGND sg13g2_buf_8
Xfanout599 _0440_ net599 VPWR VGND sg13g2_buf_8
XFILLER_46_417 VPWR VGND sg13g2_decap_4
XFILLER_25_53 VPWR VGND sg13g2_decap_8
XFILLER_42_678 VPWR VGND sg13g2_decap_4
XFILLER_10_531 VPWR VGND sg13g2_decap_4
XFILLER_2_796 VPWR VGND sg13g2_decap_8
XFILLER_38_929 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_30_clk_regs clknet_3_7__leaf_clk_regs clknet_leaf_30_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_46_995 VPWR VGND sg13g2_decap_8
XFILLER_33_612 VPWR VGND sg13g2_fill_2
XFILLER_18_686 VPWR VGND sg13g2_decap_8
XFILLER_18_697 VPWR VGND sg13g2_fill_1
X_3810_ _1700_ VPWR _0354_ VGND _1916_ net600 sg13g2_o21ai_1
X_3741_ VGND VPWR net798 _1641_ _1642_ net796 sg13g2_a21oi_1
X_3672_ VGND VPWR net807 _1990_ _1576_ net799 sg13g2_a21oi_1
X_2623_ net947 VPWR _0016_ VGND _1929_ _0835_ sg13g2_o21ai_1
X_2554_ net790 _0645_ net622 _0751_ _0781_ VPWR VGND sg13g2_or4_1
X_2485_ net752 net756 _0713_ VPWR VGND sg13g2_nor2_1
X_4224_ net669 VGND VPWR net69 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[70\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_4155_ net660 VGND VPWR net550 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[1\]
+ clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
X_3106_ _1169_ VPWR _0180_ VGND net268 _1170_ sg13g2_o21ai_1
X_4086_ _1023_ net834 _1031_ _1904_ VPWR VGND sg13g2_mux2_1
X_3037_ _1127_ net742 net638 VPWR VGND sg13g2_nand2_1
XFILLER_12_807 VPWR VGND sg13g2_fill_2
X_3939_ VGND VPWR _0910_ _1795_ _1796_ _0909_ sg13g2_a21oi_1
XFILLER_47_726 VPWR VGND sg13g2_decap_8
XFILLER_28_951 VPWR VGND sg13g2_decap_8
XFILLER_46_269 VPWR VGND sg13g2_decap_8
XFILLER_43_954 VPWR VGND sg13g2_decap_8
XFILLER_42_453 VPWR VGND sg13g2_fill_2
XFILLER_7_811 VPWR VGND sg13g2_fill_2
XFILLER_2_582 VPWR VGND sg13g2_fill_2
X_2270_ _0501_ _0492_ _0502_ VPWR VGND sg13g2_nor2b_1
XFILLER_46_781 VPWR VGND sg13g2_decap_8
XFILLER_34_987 VPWR VGND sg13g2_decap_8
XFILLER_20_158 VPWR VGND sg13g2_decap_4
X_3724_ _1613_ VPWR _1626_ VGND net795 _1625_ sg13g2_o21ai_1
X_3655_ _1559_ VPWR _1560_ VGND net796 _1554_ sg13g2_o21ai_1
X_2606_ _0825_ net588 _0824_ VPWR VGND sg13g2_nand2_1
X_3586_ _0335_ _1493_ _1967_ net583 _1956_ VPWR VGND sg13g2_a22oi_1
XFILLER_0_519 VPWR VGND sg13g2_decap_8
X_2537_ VGND VPWR _0661_ _0763_ _0764_ _0750_ sg13g2_a21oi_1
X_2468_ _0680_ VPWR _0696_ VGND _0650_ _0695_ sg13g2_o21ai_1
X_4207_ net668 VGND VPWR net241 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[53\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_2399_ VPWR VGND net742 _0629_ _0628_ net589 _0062_ _0626_ sg13g2_a221oi_1
X_4138_ net729 VGND VPWR net930 u_usb_cdc.u_sie.u_phy_rx.state_q\[3\] clknet_leaf_25_clk_regs
+ sg13g2_dfrbpq_1
X_4069_ net625 _1853_ u_usb_cdc.u_sie.u_phy_tx.data_q\[0\] _1892_ VPWR VGND _1891_
+ sg13g2_nand4_1
XFILLER_44_707 VPWR VGND sg13g2_decap_8
XFILLER_43_228 VPWR VGND sg13g2_fill_2
XFILLER_25_976 VPWR VGND sg13g2_decap_8
XFILLER_40_957 VPWR VGND sg13g2_decap_8
XFILLER_12_659 VPWR VGND sg13g2_fill_2
XFILLER_22_32 VPWR VGND sg13g2_fill_2
Xheichips25_usb_cdc_39 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_3_379 VPWR VGND sg13g2_decap_8
XFILLER_3_346 VPWR VGND sg13g2_decap_4
XFILLER_35_707 VPWR VGND sg13g2_fill_2
XFILLER_43_762 VPWR VGND sg13g2_decap_8
XFILLER_10_191 VPWR VGND sg13g2_fill_2
Xhold608 _0289_ VPWR VGND net927 sg13g2_dlygate4sd3_1
X_3440_ net566 net581 _1406_ VPWR VGND sg13g2_nor2_1
Xhold619 _0048_ VPWR VGND net938 sg13g2_dlygate4sd3_1
X_3371_ net951 _1280_ _1360_ _0254_ VPWR VGND sg13g2_mux2_1
X_2322_ net849 _0551_ _0552_ _0553_ _0554_ VPWR VGND sg13g2_nor4_1
X_2253_ _0485_ _0483_ _0484_ VPWR VGND sg13g2_xnor2_1
X_2184_ _2038_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\]
+ VPWR VGND sg13g2_nand2_2
XFILLER_26_707 VPWR VGND sg13g2_fill_1
XFILLER_38_578 VPWR VGND sg13g2_fill_1
XFILLER_25_217 VPWR VGND sg13g2_decap_4
XFILLER_19_781 VPWR VGND sg13g2_decap_4
XFILLER_34_784 VPWR VGND sg13g2_fill_2
X_3707_ VPWR VGND _1499_ net627 _1609_ net637 _1610_ _1599_ sg13g2_a221oi_1
X_3638_ net781 VPWR _1543_ VGND net785 _1441_ sg13g2_o21ai_1
X_3569_ _0877_ _1490_ _1972_ _1491_ VPWR VGND sg13g2_nand3_1
XFILLER_0_316 VPWR VGND sg13g2_decap_8
XFILLER_44_537 VPWR VGND sg13g2_fill_2
XFILLER_12_478 VPWR VGND sg13g2_decap_8
XFILLER_48_843 VPWR VGND sg13g2_decap_8
Xhold5 u_usb_cdc.u_sie.u_phy_rx.dn_q\[1\] VPWR VGND net48 sg13g2_dlygate4sd3_1
X_2940_ net515 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ _1077_ _0107_ VPWR VGND sg13g2_mux2_1
X_2871_ net9 net1020 net646 _0082_ VPWR VGND sg13g2_mux2_1
XFILLER_8_950 VPWR VGND sg13g2_decap_8
X_4472_ net733 VGND VPWR net454 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] clknet_leaf_30_clk_regs
+ sg13g2_dfrbpq_2
Xhold405 u_usb_cdc.u_sie.addr_q\[3\] VPWR VGND net448 sg13g2_dlygate4sd3_1
Xhold416 _0057_ VPWR VGND net459 sg13g2_dlygate4sd3_1
Xhold427 _0141_ VPWR VGND net470 sg13g2_dlygate4sd3_1
Xhold449 u_usb_cdc.u_ctrl_endp.class_q VPWR VGND net492 sg13g2_dlygate4sd3_1
X_3423_ net861 net428 _1397_ _0270_ VPWR VGND sg13g2_mux2_1
Xhold438 _0060_ VPWR VGND net481 sg13g2_dlygate4sd3_1
X_3354_ _1349_ VPWR _1350_ VGND _1347_ _1348_ sg13g2_o21ai_1
X_3285_ net816 net812 _1287_ VPWR VGND sg13g2_nor2_1
X_2305_ _0537_ net776 VPWR VGND net775 sg13g2_nand2b_2
X_2236_ _0468_ _0464_ _0467_ VPWR VGND sg13g2_xnor2_1
X_2167_ net717 _2022_ _2023_ VPWR VGND sg13g2_nor2_2
X_2098_ VPWR _1955_ u_usb_cdc.u_sie.crc16_q\[13\] VGND sg13g2_inv_1
XFILLER_0_1021 VPWR VGND sg13g2_decap_8
XFILLER_16_1018 VPWR VGND sg13g2_decap_8
XFILLER_1_636 VPWR VGND sg13g2_decap_8
XFILLER_0_157 VPWR VGND sg13g2_fill_1
XFILLER_49_618 VPWR VGND sg13g2_decap_8
XFILLER_13_710 VPWR VGND sg13g2_fill_1
XFILLER_12_220 VPWR VGND sg13g2_fill_2
XFILLER_40_573 VPWR VGND sg13g2_fill_2
XFILLER_5_942 VPWR VGND sg13g2_decap_8
XFILLER_4_430 VPWR VGND sg13g2_fill_2
X_3070_ _1145_ VPWR _0169_ VGND _1913_ net634 sg13g2_o21ai_1
XFILLER_39_117 VPWR VGND sg13g2_fill_2
XFILLER_48_640 VPWR VGND sg13g2_decap_8
XFILLER_16_581 VPWR VGND sg13g2_fill_2
X_3972_ net285 VPWR _0402_ VGND _1949_ net614 sg13g2_o21ai_1
X_2923_ _1065_ VPWR _0101_ VGND net618 _1066_ sg13g2_o21ai_1
XFILLER_31_540 VPWR VGND sg13g2_fill_1
X_2854_ net1044 net977 _1025_ VPWR VGND sg13g2_xor2_1
X_2785_ u_usb_cdc.u_ctrl_endp.endp_q\[1\] _1970_ net545 net500 _0962_ VPWR VGND sg13g2_nor4_1
Xhold202 _0248_ VPWR VGND net245 sg13g2_dlygate4sd3_1
Xhold213 _0173_ VPWR VGND net256 sg13g2_dlygate4sd3_1
Xhold235 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[11\] VPWR
+ VGND net278 sg13g2_dlygate4sd3_1
Xhold224 _0404_ VPWR VGND net267 sg13g2_dlygate4sd3_1
Xhold246 _0169_ VPWR VGND net289 sg13g2_dlygate4sd3_1
Xhold257 _0073_ VPWR VGND net300 sg13g2_dlygate4sd3_1
XFILLER_49_19 VPWR VGND sg13g2_decap_8
X_4455_ net726 VGND VPWR net320 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[13\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
Xhold268 _0365_ VPWR VGND net311 sg13g2_dlygate4sd3_1
X_4386_ net728 VGND VPWR net415 u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_2
X_3406_ _0611_ _0616_ _0644_ _1388_ VGND VPWR _0665_ sg13g2_nor4_2
Xfanout704 net705 net704 VPWR VGND sg13g2_buf_8
Xhold279 _0321_ VPWR VGND net322 sg13g2_dlygate4sd3_1
Xfanout715 net716 net715 VPWR VGND sg13g2_buf_8
X_3337_ _1333_ VPWR _1334_ VGND net822 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[5\]
+ sg13g2_o21ai_1
Xfanout726 net738 net726 VPWR VGND sg13g2_buf_8
Xfanout748 net749 net748 VPWR VGND sg13g2_buf_8
Xfanout737 net738 net737 VPWR VGND sg13g2_buf_8
Xfanout759 net298 net759 VPWR VGND sg13g2_buf_8
X_3268_ _1264_ net892 _1272_ _0240_ VPWR VGND sg13g2_a21o_1
X_3199_ net347 net630 _1226_ VPWR VGND sg13g2_nor2_1
X_2219_ _1932_ net944 _0451_ VPWR VGND sg13g2_nor2_2
XFILLER_42_805 VPWR VGND sg13g2_decap_4
XFILLER_42_827 VPWR VGND sg13g2_fill_2
XFILLER_41_315 VPWR VGND sg13g2_decap_4
XFILLER_10_724 VPWR VGND sg13g2_decap_4
XFILLER_10_713 VPWR VGND sg13g2_fill_2
XFILLER_6_717 VPWR VGND sg13g2_fill_1
XFILLER_10_757 VPWR VGND sg13g2_decap_8
XFILLER_2_989 VPWR VGND sg13g2_decap_8
XFILLER_39_30 VPWR VGND sg13g2_fill_2
XFILLER_49_415 VPWR VGND sg13g2_decap_8
XFILLER_39_74 VPWR VGND sg13g2_fill_1
XFILLER_18_824 VPWR VGND sg13g2_fill_1
XFILLER_45_610 VPWR VGND sg13g2_fill_1
XFILLER_45_698 VPWR VGND sg13g2_decap_8
XFILLER_13_584 VPWR VGND sg13g2_decap_4
XFILLER_9_511 VPWR VGND sg13g2_decap_8
X_2570_ _0788_ _0794_ _0700_ _0795_ VPWR VGND sg13g2_nand3_1
X_4240_ net673 VGND VPWR net289 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[2\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_4171_ net666 VGND VPWR net169 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[17\]
+ clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
X_3122_ _1182_ net761 _1141_ VPWR VGND sg13g2_nand2_2
XFILLER_49_982 VPWR VGND sg13g2_decap_8
X_3053_ _1128_ _1133_ u_usb_cdc.sie_in_data_ack _1135_ VPWR VGND sg13g2_nand3_1
XFILLER_48_492 VPWR VGND sg13g2_decap_8
X_3955_ net955 net413 _1806_ VPWR VGND sg13g2_nor2_2
XFILLER_32_860 VPWR VGND sg13g2_fill_1
X_2906_ _1053_ VPWR _0096_ VGND net619 _1054_ sg13g2_o21ai_1
X_3886_ _1755_ _1757_ _0373_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_0_clk_regs clknet_3_0__leaf_clk_regs clknet_leaf_0_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2837_ net626 _1008_ _1009_ VPWR VGND sg13g2_nor2b_1
X_2768_ _0946_ _0452_ _0450_ VPWR VGND sg13g2_nand2b_1
X_2699_ _2037_ _0884_ _2032_ _0898_ VPWR VGND sg13g2_nand3_1
X_4507_ net703 VGND VPWR net405 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[2\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_1
X_4438_ net730 VGND VPWR net339 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[5\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_1
X_4369_ net692 VGND VPWR _0297_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[2\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_47_908 VPWR VGND sg13g2_decap_8
Xfanout578 _1390_ net578 VPWR VGND sg13g2_buf_8
Xfanout589 _0622_ net589 VPWR VGND sg13g2_buf_1
XFILLER_42_613 VPWR VGND sg13g2_decap_4
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_fill_1
XFILLER_1_285 VPWR VGND sg13g2_fill_1
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_234 VPWR VGND sg13g2_fill_2
XFILLER_46_974 VPWR VGND sg13g2_decap_8
XFILLER_33_646 VPWR VGND sg13g2_fill_1
X_3740_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[21\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[29\]
+ net804 _1641_ VPWR VGND sg13g2_mux2_1
XFILLER_12_1010 VPWR VGND sg13g2_decap_8
X_3671_ net803 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[2\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[10\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[18\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[26\]
+ net799 _1575_ VPWR VGND sg13g2_mux4_1
X_2622_ net588 _0665_ net946 _0836_ VPWR VGND _0823_ sg13g2_nand4_1
X_2553_ VGND VPWR _0777_ _0779_ _0780_ _0639_ sg13g2_a21oi_1
X_2484_ _0610_ _0613_ net850 _0712_ VPWR VGND sg13g2_nand3_1
X_4223_ net669 VGND VPWR net140 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[69\]
+ clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_4154_ net680 VGND VPWR net462 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[0\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
X_3105_ net832 _1159_ u_usb_cdc.sie_out_data\[5\] _1170_ VPWR VGND sg13g2_nand3_1
X_4085_ _1903_ VPWR _0426_ VGND _1919_ _1902_ sg13g2_o21ai_1
X_3036_ _1126_ VPWR _0154_ VGND _1095_ _1098_ sg13g2_o21ai_1
XFILLER_37_985 VPWR VGND sg13g2_decap_8
XFILLER_24_602 VPWR VGND sg13g2_fill_2
XFILLER_36_484 VPWR VGND sg13g2_decap_4
XFILLER_23_123 VPWR VGND sg13g2_fill_2
XFILLER_24_668 VPWR VGND sg13g2_fill_1
X_3938_ _1795_ _2037_ _0904_ VPWR VGND sg13g2_nand2_1
X_3869_ _1978_ _2003_ _1744_ VPWR VGND sg13g2_nor2_2
XFILLER_47_705 VPWR VGND sg13g2_decap_8
XFILLER_28_930 VPWR VGND sg13g2_decap_8
XFILLER_36_53 VPWR VGND sg13g2_fill_1
XFILLER_43_933 VPWR VGND sg13g2_decap_8
XFILLER_27_484 VPWR VGND sg13g2_decap_8
XFILLER_42_410 VPWR VGND sg13g2_fill_2
XFILLER_38_738 VPWR VGND sg13g2_fill_1
XFILLER_37_248 VPWR VGND sg13g2_decap_4
XFILLER_46_760 VPWR VGND sg13g2_decap_8
XFILLER_18_484 VPWR VGND sg13g2_fill_1
XFILLER_45_281 VPWR VGND sg13g2_decap_8
XFILLER_34_966 VPWR VGND sg13g2_decap_8
XFILLER_21_605 VPWR VGND sg13g2_fill_2
XFILLER_14_690 VPWR VGND sg13g2_fill_2
XFILLER_20_137 VPWR VGND sg13g2_decap_8
X_3723_ _1618_ VPWR _1625_ VGND _1621_ _1624_ sg13g2_o21ai_1
X_3654_ _1559_ _1556_ _1558_ VPWR VGND sg13g2_nand2_1
X_2605_ net946 _0666_ _0822_ _0824_ VPWR VGND sg13g2_nor3_1
X_3585_ _0334_ net579 _1964_ net583 _1957_ VPWR VGND sg13g2_a22oi_1
X_2536_ VGND VPWR _0763_ _0762_ _0635_ sg13g2_or2_1
X_2467_ _0695_ net763 _0692_ VPWR VGND sg13g2_nand2_2
X_4206_ net662 VGND VPWR net136 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[52\]
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
X_2398_ net541 _0619_ _0629_ VPWR VGND sg13g2_nor2_1
X_4137_ net727 VGND VPWR _0034_ u_usb_cdc.u_sie.u_phy_rx.state_q\[2\] clknet_leaf_23_clk_regs
+ sg13g2_dfrbpq_1
X_4068_ _1891_ _1979_ _0434_ VPWR VGND sg13g2_nand2_1
X_3019_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ net477 _1117_ _0146_ VPWR VGND sg13g2_mux2_1
XFILLER_22_11 VPWR VGND sg13g2_fill_2
XFILLER_20_660 VPWR VGND sg13g2_decap_4
XFILLER_3_358 VPWR VGND sg13g2_decap_8
XFILLER_26_1009 VPWR VGND sg13g2_decap_8
XFILLER_47_513 VPWR VGND sg13g2_fill_2
XFILLER_35_719 VPWR VGND sg13g2_fill_2
XFILLER_28_782 VPWR VGND sg13g2_fill_2
XFILLER_27_281 VPWR VGND sg13g2_decap_4
XFILLER_43_741 VPWR VGND sg13g2_fill_1
XFILLER_15_498 VPWR VGND sg13g2_decap_4
Xhold609 u_usb_cdc.u_sie.crc16_q\[15\] VPWR VGND net928 sg13g2_dlygate4sd3_1
X_3370_ net940 _1274_ _1360_ _0253_ VPWR VGND sg13g2_mux2_1
X_2321_ u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\] u_usb_cdc.u_ctrl_endp.req_q\[4\] _0553_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_3_870 VPWR VGND sg13g2_fill_1
X_2252_ net767 u_usb_cdc.u_sie.crc16_q\[15\] _0484_ VPWR VGND sg13g2_xor2_1
XFILLER_33_4 VPWR VGND sg13g2_decap_8
X_2183_ _2037_ _1943_ _1944_ VPWR VGND sg13g2_nand2_2
XFILLER_19_760 VPWR VGND sg13g2_fill_2
XFILLER_22_914 VPWR VGND sg13g2_fill_2
X_3706_ _1600_ VPWR _1609_ VGND _1604_ _1608_ sg13g2_o21ai_1
X_3637_ _1542_ _1541_ net773 VPWR VGND sg13g2_nand2b_1
XFILLER_1_818 VPWR VGND sg13g2_fill_2
X_3568_ net842 net847 _1490_ VPWR VGND sg13g2_nor2_2
X_2519_ _0744_ _0745_ _0695_ _0746_ VPWR VGND sg13g2_nand3_1
X_3499_ VGND VPWR _1446_ _0655_ _0541_ sg13g2_or2_1
XFILLER_29_546 VPWR VGND sg13g2_fill_2
XFILLER_29_557 VPWR VGND sg13g2_decap_8
XFILLER_25_774 VPWR VGND sg13g2_decap_4
XFILLER_40_788 VPWR VGND sg13g2_fill_1
XFILLER_33_98 VPWR VGND sg13g2_fill_1
XFILLER_32_1024 VPWR VGND sg13g2_decap_4
XFILLER_48_822 VPWR VGND sg13g2_decap_8
XFILLER_0_895 VPWR VGND sg13g2_decap_8
Xhold6 u_usb_cdc.clk_cnt_q\[0\] VPWR VGND net49 sg13g2_dlygate4sd3_1
XFILLER_48_899 VPWR VGND sg13g2_decap_8
XFILLER_16_741 VPWR VGND sg13g2_decap_8
XFILLER_16_763 VPWR VGND sg13g2_fill_1
XFILLER_43_571 VPWR VGND sg13g2_fill_2
X_2870_ net8 net1010 net646 _0081_ VPWR VGND sg13g2_mux2_1
XFILLER_31_766 VPWR VGND sg13g2_fill_1
XFILLER_31_799 VPWR VGND sg13g2_fill_2
X_4471_ net736 VGND VPWR net558 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[1\] clknet_leaf_27_clk_regs
+ sg13g2_dfrbpq_2
Xhold406 u_usb_cdc.u_sie.addr_q\[1\] VPWR VGND net449 sg13g2_dlygate4sd3_1
Xhold417 _1882_ VPWR VGND net460 sg13g2_dlygate4sd3_1
X_3422_ net905 net485 _1397_ _0269_ VPWR VGND sg13g2_mux2_1
Xhold428 u_usb_cdc.u_ctrl_endp.state_q\[5\] VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold439 _0420_ VPWR VGND net482 sg13g2_dlygate4sd3_1
X_3353_ VGND VPWR _1341_ _1343_ _1349_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[3\]
+ sg13g2_a21oi_1
X_3284_ _1286_ net816 _1982_ VPWR VGND sg13g2_nand2_2
X_2304_ net790 _0535_ _0536_ VPWR VGND sg13g2_and2_1
XFILLER_39_833 VPWR VGND sg13g2_fill_2
X_2235_ _0467_ net761 net757 VPWR VGND sg13g2_xnor2_1
X_2166_ _2022_ _2021_ VPWR VGND sg13g2_inv_2
XFILLER_0_1000 VPWR VGND sg13g2_decap_8
X_2097_ VPWR _1954_ net910 VGND sg13g2_inv_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_34_582 VPWR VGND sg13g2_fill_2
XFILLER_22_733 VPWR VGND sg13g2_fill_2
XFILLER_22_766 VPWR VGND sg13g2_fill_2
X_2999_ _1111_ net253 _1108_ VPWR VGND sg13g2_nand2_1
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_45_869 VPWR VGND sg13g2_decap_8
XFILLER_44_324 VPWR VGND sg13g2_decap_4
XFILLER_44_379 VPWR VGND sg13g2_fill_2
XFILLER_13_766 VPWR VGND sg13g2_fill_1
XFILLER_8_225 VPWR VGND sg13g2_fill_1
XFILLER_8_236 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_24_clk_regs clknet_3_6__leaf_clk_regs clknet_leaf_24_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_4_453 VPWR VGND sg13g2_fill_2
XFILLER_5_998 VPWR VGND sg13g2_decap_8
XFILLER_0_692 VPWR VGND sg13g2_decap_8
XFILLER_48_696 VPWR VGND sg13g2_decap_8
X_3971_ _1814_ net284 _0942_ VPWR VGND sg13g2_nand2_1
X_2922_ _1066_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net644 VPWR VGND sg13g2_nand2_1
XFILLER_31_563 VPWR VGND sg13g2_fill_1
X_2853_ _1024_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[0\] _1023_
+ VPWR VGND sg13g2_xnor2_1
X_2784_ net850 u_usb_cdc.u_ctrl_endp.state_q\[6\] _0551_ _0747_ _0961_ VPWR VGND sg13g2_nor4_1
XFILLER_8_770 VPWR VGND sg13g2_decap_4
Xhold214 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[32\] VPWR
+ VGND net257 sg13g2_dlygate4sd3_1
Xhold203 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[38\] VPWR
+ VGND net246 sg13g2_dlygate4sd3_1
Xhold225 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[2\] VPWR
+ VGND net268 sg13g2_dlygate4sd3_1
Xhold269 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[1\] VPWR VGND net312 sg13g2_dlygate4sd3_1
Xhold247 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[26\] VPWR
+ VGND net290 sg13g2_dlygate4sd3_1
Xhold236 _0178_ VPWR VGND net279 sg13g2_dlygate4sd3_1
Xhold258 u_usb_cdc.u_sie.phy_state_q\[5\] VPWR VGND net301 sg13g2_dlygate4sd3_1
X_4454_ net726 VGND VPWR _0382_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[12\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
X_4385_ net728 VGND VPWR net956 u_usb_cdc.u_ctrl_endp.dev_state_qq\[0\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_2
X_3405_ net624 _0671_ _1387_ VPWR VGND sg13g2_nor2_1
Xfanout705 net706 net705 VPWR VGND sg13g2_buf_8
X_3336_ _1333_ net825 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[13\]
+ VPWR VGND sg13g2_nand2b_1
Xfanout716 _1939_ net716 VPWR VGND sg13g2_buf_8
Xfanout738 net1048 net738 VPWR VGND sg13g2_buf_8
Xfanout749 u_usb_cdc.clk_gate_q net749 VPWR VGND sg13g2_buf_8
Xfanout727 net728 net727 VPWR VGND sg13g2_buf_8
X_3267_ VGND VPWR _1270_ _1271_ _1272_ _1264_ sg13g2_a21oi_1
XFILLER_22_1023 VPWR VGND sg13g2_decap_4
XFILLER_39_652 VPWR VGND sg13g2_fill_1
X_2218_ _0443_ _0445_ _0442_ _0450_ VPWR VGND _0449_ sg13g2_nand4_1
X_3198_ VGND VPWR _1913_ net630 _0217_ _1225_ sg13g2_a21oi_1
XFILLER_39_674 VPWR VGND sg13g2_decap_8
X_2149_ VPWR _2005_ net938 VGND sg13g2_inv_1
XFILLER_22_574 VPWR VGND sg13g2_fill_2
XFILLER_6_707 VPWR VGND sg13g2_fill_1
XFILLER_30_11 VPWR VGND sg13g2_fill_2
XFILLER_2_913 VPWR VGND sg13g2_decap_8
XFILLER_1_434 VPWR VGND sg13g2_fill_2
XFILLER_1_423 VPWR VGND sg13g2_decap_8
XFILLER_2_968 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_9_501 VPWR VGND sg13g2_fill_2
XFILLER_9_545 VPWR VGND sg13g2_fill_2
XFILLER_45_1023 VPWR VGND sg13g2_decap_4
X_4170_ net667 VGND VPWR net251 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[16\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_3121_ net325 net632 _1181_ VPWR VGND sg13g2_nor2_1
XFILLER_49_961 VPWR VGND sg13g2_decap_8
X_3052_ _1134_ net1037 _1133_ VPWR VGND sg13g2_nand2_1
XFILLER_48_471 VPWR VGND sg13g2_decap_8
XFILLER_35_110 VPWR VGND sg13g2_fill_1
XFILLER_17_880 VPWR VGND sg13g2_fill_1
X_3954_ VGND VPWR net747 net306 _0393_ _1805_ sg13g2_a21oi_1
X_2905_ _1054_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net645 VPWR VGND sg13g2_nand2_1
X_3885_ _1757_ _1756_ net982 VPWR VGND sg13g2_nand2b_1
X_2836_ net835 _0926_ _1008_ VPWR VGND sg13g2_nor2_2
X_2767_ u_usb_cdc.bus_reset net726 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.rstn VPWR
+ VGND sg13g2_nor2b_2
X_2698_ _0896_ VPWR _0002_ VGND _0720_ _0897_ sg13g2_o21ai_1
X_4506_ net703 VGND VPWR net390 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[1\] clknet_leaf_30_clk_regs
+ sg13g2_dfrbpq_2
X_4437_ net731 VGND VPWR net311 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[4\] clknet_leaf_26_clk_regs
+ sg13g2_dfrbpq_1
X_4368_ net692 VGND VPWR _0296_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[1\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_4299_ net673 VGND VPWR net324 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[61\]
+ clknet_leaf_47_clk_regs sg13g2_dfrbpq_1
X_3319_ VGND VPWR net818 _1997_ _1318_ net815 sg13g2_a21oi_1
Xfanout579 net580 net579 VPWR VGND sg13g2_buf_8
XFILLER_39_493 VPWR VGND sg13g2_fill_1
XFILLER_39_482 VPWR VGND sg13g2_fill_2
XFILLER_15_806 VPWR VGND sg13g2_fill_2
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_6_526 VPWR VGND sg13g2_fill_2
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_6_537 VPWR VGND sg13g2_fill_2
XFILLER_1_297 VPWR VGND sg13g2_decap_8
XFILLER_2_59 VPWR VGND sg13g2_fill_2
XFILLER_18_611 VPWR VGND sg13g2_decap_4
XFILLER_46_953 VPWR VGND sg13g2_decap_8
XFILLER_45_430 VPWR VGND sg13g2_decap_8
XFILLER_17_143 VPWR VGND sg13g2_fill_2
XFILLER_18_666 VPWR VGND sg13g2_decap_8
XFILLER_45_463 VPWR VGND sg13g2_fill_1
XFILLER_17_176 VPWR VGND sg13g2_fill_2
X_3670_ _1574_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[66\] net628
+ VPWR VGND sg13g2_nand2_1
X_2621_ VPWR VGND _0610_ net591 _0834_ _0549_ _0835_ net589 sg13g2_a221oi_1
X_2552_ _0779_ _0698_ _0778_ u_usb_cdc.u_ctrl_endp.req_q\[7\] net757 VPWR VGND sg13g2_a22oi_1
X_2483_ net763 net762 _0708_ _0710_ _0711_ VPWR VGND sg13g2_or4_1
X_4222_ net669 VGND VPWR net134 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[68\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
X_4153_ net663 VGND VPWR _0082_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_2
X_3104_ _1169_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[13\]
+ _1151_ VPWR VGND sg13g2_nand2_1
X_4084_ _1903_ net164 _1902_ VPWR VGND sg13g2_nand2_1
X_3035_ _1126_ net137 _1118_ VPWR VGND sg13g2_nand2_1
XFILLER_23_146 VPWR VGND sg13g2_decap_8
X_3937_ _0387_ _1794_ _1976_ _1793_ _0916_ VPWR VGND sg13g2_a22oi_1
XFILLER_32_680 VPWR VGND sg13g2_fill_1
X_3868_ VGND VPWR _0369_ _1743_ _1742_ sg13g2_or2_1
XFILLER_20_886 VPWR VGND sg13g2_fill_2
X_3799_ net592 _1692_ net765 _1695_ VPWR VGND sg13g2_nand3_1
X_2819_ _0962_ u_usb_cdc.u_ctrl_endp.in_endp_q net851 _0994_ VPWR VGND sg13g2_a21o_1
XFILLER_4_1009 VPWR VGND sg13g2_decap_8
XFILLER_43_912 VPWR VGND sg13g2_decap_8
XFILLER_15_603 VPWR VGND sg13g2_fill_2
XFILLER_28_986 VPWR VGND sg13g2_decap_8
XFILLER_14_113 VPWR VGND sg13g2_fill_1
XFILLER_14_124 VPWR VGND sg13g2_fill_2
XFILLER_43_989 VPWR VGND sg13g2_decap_8
XFILLER_35_1011 VPWR VGND sg13g2_decap_8
XFILLER_10_341 VPWR VGND sg13g2_decap_4
XFILLER_10_396 VPWR VGND sg13g2_fill_1
XFILLER_42_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_127 VPWR VGND sg13g2_fill_1
X_3722_ net796 VPWR _1624_ VGND _1622_ _1623_ sg13g2_o21ai_1
X_3653_ VGND VPWR net802 _1557_ _1558_ _1923_ sg13g2_a21oi_1
X_2604_ VPWR _0823_ _0822_ VGND sg13g2_inv_1
XFILLER_6_890 VPWR VGND sg13g2_fill_1
X_3584_ _0333_ net580 _1965_ net583 _1958_ VPWR VGND sg13g2_a22oi_1
X_2535_ _0761_ VPWR _0762_ VGND net784 _0540_ sg13g2_o21ai_1
X_2466_ net723 _0693_ _0694_ VPWR VGND sg13g2_nor2_1
X_4205_ net660 VGND VPWR net87 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[51\]
+ clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
X_2397_ VGND VPWR _0607_ _0627_ _0628_ _0612_ sg13g2_a21oi_1
X_4136_ net727 VGND VPWR net395 u_usb_cdc.u_sie.u_phy_rx.state_q\[1\] clknet_leaf_25_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_238 VPWR VGND sg13g2_decap_4
X_4067_ _1890_ VPWR _0421_ VGND net748 _2003_ sg13g2_o21ai_1
X_3018_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ net479 _1117_ _0145_ VPWR VGND sg13g2_mux2_1
XFILLER_11_105 VPWR VGND sg13g2_fill_2
XFILLER_3_304 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_49_clk_regs clknet_3_1__leaf_clk_regs clknet_leaf_49_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_16_901 VPWR VGND sg13g2_decap_4
XFILLER_35_709 VPWR VGND sg13g2_fill_1
XFILLER_16_934 VPWR VGND sg13g2_fill_2
XFILLER_11_683 VPWR VGND sg13g2_fill_1
XFILLER_10_193 VPWR VGND sg13g2_fill_1
X_2320_ VGND VPWR _0552_ net850 u_usb_cdc.u_ctrl_endp.state_q\[1\] sg13g2_or2_1
X_2251_ net766 u_usb_cdc.u_sie.crc16_q\[14\] _0483_ VPWR VGND sg13g2_xor2_1
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_2182_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[2\] u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\]
+ _2036_ VPWR VGND sg13g2_nor2_2
XFILLER_19_750 VPWR VGND sg13g2_fill_1
XFILLER_38_569 VPWR VGND sg13g2_decap_8
XFILLER_34_786 VPWR VGND sg13g2_fill_1
X_3705_ _1606_ VPWR _1608_ VGND net773 _1607_ sg13g2_o21ai_1
X_3636_ _0762_ _1540_ _0656_ _1541_ VPWR VGND sg13g2_nand3_1
X_3567_ _1488_ VPWR _0322_ VGND _0867_ _1489_ sg13g2_o21ai_1
X_2518_ VGND VPWR _0745_ _0727_ _0691_ sg13g2_or2_1
X_3498_ _1445_ net781 _1437_ VPWR VGND sg13g2_nand2_1
X_2449_ _0651_ _0664_ _0642_ _0679_ VPWR VGND _0677_ sg13g2_nand4_1
X_4119_ net699 VGND VPWR _0020_ u_usb_cdc.u_sie.phy_state_q\[1\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_44_539 VPWR VGND sg13g2_fill_1
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_40_734 VPWR VGND sg13g2_fill_2
XFILLER_32_1003 VPWR VGND sg13g2_decap_8
XFILLER_4_668 VPWR VGND sg13g2_fill_1
XFILLER_48_801 VPWR VGND sg13g2_decap_8
XFILLER_0_874 VPWR VGND sg13g2_decap_8
Xhold7 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[68\] VPWR VGND
+ net50 sg13g2_dlygate4sd3_1
XFILLER_48_878 VPWR VGND sg13g2_decap_8
X_4470_ net736 VGND VPWR net555 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[0\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_8_985 VPWR VGND sg13g2_decap_8
Xhold418 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[0\] VPWR VGND
+ net461 sg13g2_dlygate4sd3_1
Xhold407 u_usb_cdc.u_sie.u_phy_rx.rx_valid_q VPWR VGND net450 sg13g2_dlygate4sd3_1
X_3421_ net868 net499 _1397_ _0268_ VPWR VGND sg13g2_mux2_1
Xhold429 _0015_ VPWR VGND net472 sg13g2_dlygate4sd3_1
X_3352_ net813 VPWR _1348_ VGND net814 _1345_ sg13g2_o21ai_1
X_2303_ net791 net787 net779 _0535_ VPWR VGND sg13g2_nor3_1
X_3283_ net824 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[32\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[40\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[48\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[56\] net816 _1285_
+ VPWR VGND sg13g2_mux4_1
XFILLER_39_845 VPWR VGND sg13g2_fill_2
X_2234_ _0466_ _0461_ _0465_ VPWR VGND sg13g2_xnor2_1
X_2165_ u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[1\] u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[2\]
+ _2021_ VPWR VGND u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] sg13g2_nand3b_1
XFILLER_0_70 VPWR VGND sg13g2_decap_8
X_2096_ VPWR _1953_ net928 VGND sg13g2_inv_1
X_2998_ _1110_ VPWR _0132_ VGND _1064_ net610 sg13g2_o21ai_1
X_3619_ _1525_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[64\] net628
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_44_314 VPWR VGND sg13g2_fill_1
XFILLER_45_848 VPWR VGND sg13g2_decap_8
XFILLER_12_222 VPWR VGND sg13g2_fill_1
XFILLER_40_542 VPWR VGND sg13g2_fill_2
XFILLER_5_911 VPWR VGND sg13g2_decap_4
XFILLER_4_432 VPWR VGND sg13g2_fill_1
XFILLER_5_977 VPWR VGND sg13g2_decap_8
XFILLER_0_671 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_fill_1
XFILLER_48_675 VPWR VGND sg13g2_decap_8
XFILLER_39_1009 VPWR VGND sg13g2_decap_8
X_3970_ _1813_ VPWR _0401_ VGND _1947_ net614 sg13g2_o21ai_1
XFILLER_16_594 VPWR VGND sg13g2_fill_2
XFILLER_16_583 VPWR VGND sg13g2_fill_1
X_2921_ _1065_ net182 _1060_ VPWR VGND sg13g2_nand2_1
X_2852_ VGND VPWR net834 _1023_ _1019_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ sg13g2_a21oi_2
X_2783_ _0958_ _0959_ _0960_ _0067_ VPWR VGND sg13g2_nor3_1
Xhold204 _0205_ VPWR VGND net247 sg13g2_dlygate4sd3_1
Xhold215 _0199_ VPWR VGND net258 sg13g2_dlygate4sd3_1
Xhold226 _0180_ VPWR VGND net269 sg13g2_dlygate4sd3_1
X_4453_ net726 VGND VPWR net438 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[11\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_2
Xhold248 _0193_ VPWR VGND net291 sg13g2_dlygate4sd3_1
Xhold237 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[28\] VPWR
+ VGND net280 sg13g2_dlygate4sd3_1
Xhold259 _0024_ VPWR VGND net302 sg13g2_dlygate4sd3_1
X_3404_ _1386_ net980 _1369_ _0262_ VPWR VGND sg13g2_mux2_1
X_4384_ net677 VGND VPWR net410 u_usb_cdc.u_sie.addr_q\[6\] clknet_leaf_49_clk_regs
+ sg13g2_dfrbpq_1
Xfanout706 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.rstn net706 VPWR VGND sg13g2_buf_8
X_3335_ net821 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[37\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[45\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[53\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[61\] net816 _1332_
+ VPWR VGND sg13g2_mux4_1
Xfanout739 net741 net739 VPWR VGND sg13g2_buf_8
Xfanout717 _1939_ net717 VPWR VGND sg13g2_buf_8
Xfanout728 net738 net728 VPWR VGND sg13g2_buf_8
X_3266_ _1271_ _0604_ _1269_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[1\]
+ net755 VPWR VGND sg13g2_a22oi_1
X_2217_ _0444_ _0446_ _0447_ _0448_ _0449_ VPWR VGND sg13g2_nor4_1
X_3197_ net416 net630 _1225_ VPWR VGND sg13g2_nor2_1
X_2148_ VPWR _2004_ net387 VGND sg13g2_inv_1
X_2079_ VPWR _1936_ u_usb_cdc.u_ctrl_endp.rec_q\[0\] VGND sg13g2_inv_1
XFILLER_22_553 VPWR VGND sg13g2_fill_2
XFILLER_1_402 VPWR VGND sg13g2_decap_8
XFILLER_2_947 VPWR VGND sg13g2_decap_8
XFILLER_1_468 VPWR VGND sg13g2_fill_2
XFILLER_7_1007 VPWR VGND sg13g2_decap_8
XFILLER_39_32 VPWR VGND sg13g2_fill_1
XFILLER_44_144 VPWR VGND sg13g2_fill_2
XFILLER_9_568 VPWR VGND sg13g2_fill_2
XFILLER_9_579 VPWR VGND sg13g2_fill_1
XFILLER_45_1002 VPWR VGND sg13g2_decap_8
X_3120_ VGND VPWR _1176_ _1180_ _0184_ net441 sg13g2_a21oi_1
XFILLER_49_940 VPWR VGND sg13g2_decap_8
X_3051_ _1133_ net1034 net639 VPWR VGND sg13g2_nand2_2
XFILLER_48_450 VPWR VGND sg13g2_decap_8
XFILLER_36_601 VPWR VGND sg13g2_fill_2
XFILLER_36_667 VPWR VGND sg13g2_fill_2
X_3953_ net754 net747 _1805_ VPWR VGND sg13g2_nor2_1
XFILLER_32_840 VPWR VGND sg13g2_fill_2
XFILLER_35_199 VPWR VGND sg13g2_fill_1
X_2904_ _1053_ net131 _1037_ VPWR VGND sg13g2_nand2_1
X_3884_ net361 net365 net741 _1756_ VPWR VGND net336 sg13g2_nand4_1
X_2835_ _1007_ net299 net718 VPWR VGND sg13g2_nand2_1
X_2766_ net49 net61 _0040_ VPWR VGND sg13g2_xor2_1
X_2697_ net623 _0706_ net794 _0897_ VPWR VGND sg13g2_nand3_1
X_4505_ net703 VGND VPWR net351 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[0\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
X_4436_ net730 VGND VPWR net330 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_2
X_4367_ net692 VGND VPWR _0295_ u_usb_cdc.u_ctrl_endp.byte_cnt_q\[0\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
X_3318_ VGND VPWR net815 _1316_ _1317_ net812 sg13g2_a21oi_1
X_4298_ net672 VGND VPWR _0227_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[60\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_3249_ _1254_ net814 _1255_ VPWR VGND sg13g2_xor2_1
XFILLER_26_177 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_fill_1
XFILLER_41_136 VPWR VGND sg13g2_fill_2
XFILLER_42_659 VPWR VGND sg13g2_fill_2
XFILLER_2_733 VPWR VGND sg13g2_decap_8
XFILLER_29_1008 VPWR VGND sg13g2_decap_8
XFILLER_2_744 VPWR VGND sg13g2_fill_2
Xhold590 _0293_ VPWR VGND net909 sg13g2_dlygate4sd3_1
XFILLER_49_203 VPWR VGND sg13g2_fill_2
XFILLER_49_214 VPWR VGND sg13g2_fill_1
XFILLER_46_932 VPWR VGND sg13g2_decap_8
XFILLER_18_634 VPWR VGND sg13g2_decap_4
XFILLER_17_133 VPWR VGND sg13g2_fill_2
XFILLER_41_692 VPWR VGND sg13g2_fill_2
X_2620_ u_usb_cdc.sie_in_data_ack _0549_ _0595_ _0615_ _0834_ VPWR VGND sg13g2_nor4_1
X_2551_ u_usb_cdc.u_ctrl_endp.req_q\[1\] u_usb_cdc.u_ctrl_endp.req_q\[9\] _0749_ _0778_
+ VPWR VGND sg13g2_or3_1
X_2482_ _0710_ net794 _0709_ VPWR VGND sg13g2_nand2_1
X_4221_ net669 VGND VPWR net124 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[67\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
X_4152_ net663 VGND VPWR _0081_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[6\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_2
X_3103_ _1167_ VPWR _0179_ VGND net828 _1168_ sg13g2_o21ai_1
X_4083_ _1902_ net640 _1899_ VPWR VGND sg13g2_nand2_1
X_3034_ _1125_ VPWR _0153_ VGND _1093_ _1098_ sg13g2_o21ai_1
XFILLER_24_659 VPWR VGND sg13g2_fill_1
X_3936_ _1746_ _1789_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[16\] _1794_ VPWR VGND sg13g2_nand3_1
X_3867_ VPWR VGND net1007 _2039_ _0898_ _2044_ _1743_ _0881_ sg13g2_a221oi_1
X_3798_ _1694_ VPWR _0348_ VGND net721 net600 sg13g2_o21ai_1
X_2818_ _0993_ _0992_ _0566_ _0989_ net856 VPWR VGND sg13g2_a22oi_1
X_2749_ _0937_ net543 net11 VPWR VGND sg13g2_nand2b_1
X_4419_ net687 VGND VPWR _0347_ u_usb_cdc.sie_out_data\[0\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_965 VPWR VGND sg13g2_decap_8
XFILLER_36_33 VPWR VGND sg13g2_fill_1
XFILLER_39_291 VPWR VGND sg13g2_fill_2
XFILLER_42_401 VPWR VGND sg13g2_decap_4
XFILLER_42_412 VPWR VGND sg13g2_fill_1
XFILLER_43_968 VPWR VGND sg13g2_decap_8
XFILLER_7_858 VPWR VGND sg13g2_decap_8
XFILLER_2_541 VPWR VGND sg13g2_decap_8
XFILLER_34_902 VPWR VGND sg13g2_decap_4
XFILLER_46_795 VPWR VGND sg13g2_decap_8
X_3721_ net798 VPWR _1623_ VGND net805 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[52\]
+ sg13g2_o21ai_1
X_3652_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[49\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[57\]
+ net807 _1557_ VPWR VGND sg13g2_mux2_1
X_3583_ _0332_ net580 _0499_ net584 _1959_ VPWR VGND sg13g2_a22oi_1
X_2603_ net772 net942 _0546_ _0821_ _0822_ VPWR VGND sg13g2_or4_1
X_2534_ _0761_ net787 _0675_ VPWR VGND sg13g2_nand2_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_2465_ _0682_ _0689_ net721 _0693_ VPWR VGND sg13g2_nand3_1
X_4204_ net666 VGND VPWR net254 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[50\]
+ clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
X_2396_ _0550_ _0552_ _0627_ VPWR VGND sg13g2_nor2_1
XFILLER_29_729 VPWR VGND sg13g2_fill_1
X_4135_ net727 VGND VPWR _0065_ _0052_ clknet_leaf_23_clk_regs sg13g2_dfrbpq_1
XFILLER_3_1010 VPWR VGND sg13g2_decap_8
X_4066_ _2036_ _0882_ net748 _1890_ VPWR VGND sg13g2_nand3_1
X_3017_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ net463 _1117_ _0144_ VPWR VGND sg13g2_mux2_1
XFILLER_37_762 VPWR VGND sg13g2_fill_1
XFILLER_19_1018 VPWR VGND sg13g2_decap_8
XFILLER_12_618 VPWR VGND sg13g2_decap_4
XFILLER_22_13 VPWR VGND sg13g2_fill_1
X_3919_ net896 net713 _1781_ _0382_ VPWR VGND sg13g2_a21o_1
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_28_773 VPWR VGND sg13g2_fill_2
XFILLER_28_784 VPWR VGND sg13g2_fill_1
XFILLER_31_905 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_18_clk_regs clknet_3_3__leaf_clk_regs clknet_leaf_18_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_7_666 VPWR VGND sg13g2_fill_2
XFILLER_7_655 VPWR VGND sg13g2_fill_2
XFILLER_2_393 VPWR VGND sg13g2_decap_8
X_2250_ _0482_ _0480_ _0441_ VPWR VGND sg13g2_nand2b_1
X_2181_ _2034_ VPWR _2035_ VGND _1943_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[0\] sg13g2_o21ai_1
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_19_740 VPWR VGND sg13g2_fill_2
XFILLER_18_261 VPWR VGND sg13g2_fill_1
XFILLER_22_916 VPWR VGND sg13g2_fill_1
X_3704_ VGND VPWR _1607_ _0685_ net780 sg13g2_or2_1
XFILLER_30_982 VPWR VGND sg13g2_decap_8
X_3635_ _1538_ net780 _1540_ VPWR VGND sg13g2_xor2_1
X_3566_ _0584_ net400 _1489_ VPWR VGND sg13g2_xor2_1
X_2517_ _1942_ _0636_ _0744_ VPWR VGND sg13g2_nor2_1
X_3497_ _1443_ VPWR _0297_ VGND _1439_ _1444_ sg13g2_o21ai_1
X_2448_ _0664_ _0677_ _0651_ _0678_ VPWR VGND sg13g2_nand3_1
XFILLER_25_1011 VPWR VGND sg13g2_decap_8
X_2379_ _0598_ _0609_ _0610_ VPWR VGND sg13g2_nor2b_2
X_4118_ net695 VGND VPWR _0063_ _0050_ clknet_leaf_39_clk_regs sg13g2_dfrbpq_1
XFILLER_29_548 VPWR VGND sg13g2_fill_1
X_4049_ _1877_ net848 _1712_ VPWR VGND sg13g2_nand2_1
XFILLER_17_57 VPWR VGND sg13g2_decap_8
XFILLER_13_905 VPWR VGND sg13g2_decap_8
XFILLER_33_34 VPWR VGND sg13g2_decap_4
XFILLER_4_658 VPWR VGND sg13g2_decap_4
Xhold8 _1331_ VPWR VGND net51 sg13g2_dlygate4sd3_1
XFILLER_48_857 VPWR VGND sg13g2_decap_8
XFILLER_15_242 VPWR VGND sg13g2_fill_2
XFILLER_43_573 VPWR VGND sg13g2_fill_1
XFILLER_8_964 VPWR VGND sg13g2_decap_8
Xhold408 _0045_ VPWR VGND net451 sg13g2_dlygate4sd3_1
XFILLER_48_1011 VPWR VGND sg13g2_decap_8
Xhold419 _0083_ VPWR VGND net462 sg13g2_dlygate4sd3_1
X_3420_ _0588_ _0623_ _1396_ _1397_ VPWR VGND sg13g2_nor3_2
X_3351_ VGND VPWR net821 _2001_ _1347_ _1346_ sg13g2_a21oi_1
X_2302_ _0534_ net788 net793 VPWR VGND sg13g2_nand2b_1
X_3282_ _1284_ _0937_ _0936_ VPWR VGND sg13g2_nand2b_1
X_2233_ _0464_ net766 _0465_ VPWR VGND sg13g2_xor2_1
X_2164_ VGND VPWR net754 _2020_ _2019_ _2018_ sg13g2_a21oi_2
X_2095_ _1952_ net338 VPWR VGND sg13g2_inv_2
XFILLER_34_584 VPWR VGND sg13g2_fill_1
X_2997_ _1110_ net80 _1108_ VPWR VGND sg13g2_nand2_1
X_3618_ VGND VPWR _1524_ _1490_ net753 sg13g2_or2_1
X_3549_ _1478_ net354 _1476_ VPWR VGND sg13g2_nand2_1
XFILLER_12_201 VPWR VGND sg13g2_fill_1
XFILLER_44_99 VPWR VGND sg13g2_fill_2
XFILLER_8_238 VPWR VGND sg13g2_fill_1
XFILLER_5_956 VPWR VGND sg13g2_decap_8
XFILLER_4_455 VPWR VGND sg13g2_fill_1
XFILLER_0_650 VPWR VGND sg13g2_decap_8
XFILLER_47_131 VPWR VGND sg13g2_fill_1
XFILLER_48_654 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_33_clk_regs clknet_3_4__leaf_clk_regs clknet_leaf_33_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_16_551 VPWR VGND sg13g2_fill_2
XFILLER_44_893 VPWR VGND sg13g2_decap_8
X_2920_ _1063_ VPWR _0100_ VGND net618 _1064_ sg13g2_o21ai_1
XFILLER_15_1010 VPWR VGND sg13g2_decap_8
X_2851_ _1021_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[3\] _1022_
+ VPWR VGND sg13g2_xor2_1
X_2782_ net768 _1987_ _0952_ _0956_ _0960_ VPWR VGND sg13g2_nor4_1
Xhold216 net21 VPWR VGND net259 sg13g2_dlygate4sd3_1
Xhold205 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[19\] VPWR VGND
+ net248 sg13g2_dlygate4sd3_1
X_4452_ net726 VGND VPWR net341 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[10\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
Xhold238 _0195_ VPWR VGND net281 sg13g2_dlygate4sd3_1
Xhold249 u_usb_cdc.u_sie.u_phy_tx.data_q\[4\] VPWR VGND net292 sg13g2_dlygate4sd3_1
Xhold227 u_usb_cdc.u_sie.rx_data\[7\] VPWR VGND net270 sg13g2_dlygate4sd3_1
X_3403_ _1384_ VPWR _1386_ VGND _1372_ _1385_ sg13g2_o21ai_1
X_4383_ net677 VGND VPWR net382 u_usb_cdc.u_sie.addr_q\[5\] clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_1
X_3334_ VGND VPWR _2010_ net616 _0247_ net51 sg13g2_a21oi_1
Xfanout718 _1939_ net718 VPWR VGND sg13g2_buf_1
Xfanout707 net708 net707 VPWR VGND sg13g2_buf_8
Xfanout729 net731 net729 VPWR VGND sg13g2_buf_8
X_3265_ _1153_ _1193_ _0714_ _1270_ VPWR VGND sg13g2_nand3_1
X_2216_ u_usb_cdc.addr\[5\] u_usb_cdc.sie_out_data\[5\] _0448_ VPWR VGND sg13g2_xor2_1
XFILLER_39_632 VPWR VGND sg13g2_fill_1
X_3196_ VGND VPWR net722 net631 _0216_ net343 sg13g2_a21oi_1
X_2147_ VPWR _2003_ net374 VGND sg13g2_inv_1
X_2078_ VPWR _1935_ net1028 VGND sg13g2_inv_1
XFILLER_22_543 VPWR VGND sg13g2_fill_1
XFILLER_22_576 VPWR VGND sg13g2_fill_1
XFILLER_1_447 VPWR VGND sg13g2_decap_8
XFILLER_39_11 VPWR VGND sg13g2_decap_4
XFILLER_49_429 VPWR VGND sg13g2_decap_8
XFILLER_45_635 VPWR VGND sg13g2_fill_1
XFILLER_45_668 VPWR VGND sg13g2_fill_1
XFILLER_45_657 VPWR VGND sg13g2_decap_8
XFILLER_0_491 VPWR VGND sg13g2_decap_8
X_3050_ _1021_ net994 _1032_ _0162_ VPWR VGND sg13g2_mux2_1
XFILLER_49_996 VPWR VGND sg13g2_decap_8
XFILLER_35_101 VPWR VGND sg13g2_fill_2
XFILLER_36_624 VPWR VGND sg13g2_fill_2
XFILLER_36_646 VPWR VGND sg13g2_decap_8
XFILLER_17_860 VPWR VGND sg13g2_fill_2
XFILLER_17_871 VPWR VGND sg13g2_decap_8
X_3952_ VGND VPWR net747 _0945_ _0392_ _1804_ sg13g2_a21oi_1
X_2903_ _1051_ VPWR _0095_ VGND net619 _1052_ sg13g2_o21ai_1
X_3883_ net741 VPWR _1755_ VGND _1745_ _1754_ sg13g2_o21ai_1
X_2834_ VGND VPWR _1004_ _1005_ _0072_ net262 sg13g2_a21oi_1
X_2765_ VGND VPWR u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[3\] _1993_ net30 _0054_ sg13g2_a21oi_1
X_4504_ net730 VGND VPWR net375 u_usb_cdc.u_sie.u_phy_rx.se0_q clknet_leaf_26_clk_regs
+ sg13g2_dfrbpq_1
X_2696_ net894 VPWR _0896_ VGND _0812_ _0895_ sg13g2_o21ai_1
XFILLER_6_70 VPWR VGND sg13g2_fill_1
X_4435_ net730 VGND VPWR net422 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[2\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_1
X_4366_ net692 VGND VPWR net565 u_usb_cdc.u_ctrl_endp.max_length_q\[6\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_3317_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[19\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[27\]
+ net818 _1316_ VPWR VGND sg13g2_mux2_1
X_4297_ net673 VGND VPWR _0226_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[59\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_3248_ _1254_ _1153_ _1193_ VPWR VGND sg13g2_nand2_1
X_3179_ _1215_ VPWR _0208_ VGND net712 _1162_ sg13g2_o21ai_1
XFILLER_39_484 VPWR VGND sg13g2_fill_1
XFILLER_15_808 VPWR VGND sg13g2_fill_1
XFILLER_42_627 VPWR VGND sg13g2_decap_4
XFILLER_25_46 VPWR VGND sg13g2_decap_8
XFILLER_10_524 VPWR VGND sg13g2_decap_8
XFILLER_6_539 VPWR VGND sg13g2_fill_1
XFILLER_2_712 VPWR VGND sg13g2_decap_8
Xhold580 _0291_ VPWR VGND net899 sg13g2_dlygate4sd3_1
XFILLER_2_789 VPWR VGND sg13g2_decap_8
Xhold591 u_usb_cdc.u_sie.crc16_q\[14\] VPWR VGND net910 sg13g2_dlygate4sd3_1
XFILLER_2_39 VPWR VGND sg13g2_decap_4
XFILLER_46_911 VPWR VGND sg13g2_decap_8
XFILLER_18_602 VPWR VGND sg13g2_fill_2
XFILLER_17_145 VPWR VGND sg13g2_fill_1
XFILLER_46_988 VPWR VGND sg13g2_decap_8
XFILLER_17_178 VPWR VGND sg13g2_fill_1
XFILLER_12_1024 VPWR VGND sg13g2_decap_4
X_2550_ u_usb_cdc.u_ctrl_endp.req_q\[6\] VPWR _0777_ VGND _0698_ _0767_ sg13g2_o21ai_1
X_2481_ net880 net953 _0709_ VPWR VGND sg13g2_nor2_1
X_4220_ net667 VGND VPWR net110 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[66\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
X_4151_ net663 VGND VPWR _0080_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[5\]
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_2
X_3102_ net832 _1159_ net759 _1168_ VPWR VGND sg13g2_nand3_1
X_4082_ _1901_ VPWR _0425_ VGND _1919_ _1900_ sg13g2_o21ai_1
XFILLER_49_793 VPWR VGND sg13g2_decap_8
X_3033_ _1125_ net68 _1118_ VPWR VGND sg13g2_nand2_1
XFILLER_37_999 VPWR VGND sg13g2_decap_8
X_3935_ VGND VPWR _1791_ _1793_ _0386_ _1792_ sg13g2_a21oi_1
XFILLER_32_671 VPWR VGND sg13g2_decap_8
X_3866_ _0901_ net1039 _1742_ VPWR VGND sg13g2_nor2b_1
X_3797_ net592 _1692_ net766 _1694_ VPWR VGND sg13g2_nand3_1
X_2817_ u_usb_cdc.endp\[2\] _0988_ _0990_ _0991_ _0992_ VPWR VGND sg13g2_nor4_1
XFILLER_20_888 VPWR VGND sg13g2_fill_1
XFILLER_11_26 VPWR VGND sg13g2_fill_2
X_2748_ net739 VPWR _0936_ VGND _0934_ _0935_ sg13g2_o21ai_1
X_2679_ _0880_ VPWR _0019_ VGND _1920_ net601 sg13g2_o21ai_1
X_4418_ net705 VGND VPWR _0346_ u_usb_cdc.u_sie.data_q\[7\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_2
X_4349_ net676 VGND VPWR net429 u_usb_cdc.u_ctrl_endp.addr_dd\[2\] clknet_leaf_47_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_47_719 VPWR VGND sg13g2_decap_8
XFILLER_28_944 VPWR VGND sg13g2_decap_8
XFILLER_15_605 VPWR VGND sg13g2_fill_1
XFILLER_43_947 VPWR VGND sg13g2_decap_8
XFILLER_7_804 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_38_708 VPWR VGND sg13g2_fill_1
XFILLER_46_774 VPWR VGND sg13g2_decap_8
XFILLER_42_980 VPWR VGND sg13g2_decap_8
X_3720_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[60\] net805 _1622_
+ VPWR VGND sg13g2_nor2b_1
X_3651_ _1555_ VPWR _1556_ VGND net807 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[33\]
+ sg13g2_o21ai_1
X_3582_ _0331_ net580 _0498_ net584 _1961_ VPWR VGND sg13g2_a22oi_1
X_2602_ _0821_ net779 _0685_ VPWR VGND sg13g2_nand2_1
X_2533_ _0712_ _0759_ _0760_ VPWR VGND sg13g2_nor2_1
X_2464_ net762 _0691_ _0692_ VPWR VGND sg13g2_nor2_2
X_4203_ net666 VGND VPWR net81 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[49\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_2395_ net541 _0625_ _0626_ VPWR VGND net849 sg13g2_nand3b_1
X_4134_ net735 VGND VPWR net315 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[4\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_3_71 VPWR VGND sg13g2_fill_2
X_4065_ VGND VPWR _1908_ net643 _0420_ _1889_ sg13g2_a21oi_1
XFILLER_49_590 VPWR VGND sg13g2_decap_8
X_3016_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net475 _1117_ _0143_ VPWR VGND sg13g2_mux2_1
XFILLER_25_969 VPWR VGND sg13g2_decap_8
XFILLER_33_991 VPWR VGND sg13g2_decap_8
X_3918_ _1747_ _1779_ _1780_ _1781_ VPWR VGND sg13g2_nor3_1
X_3849_ _1731_ VPWR _0362_ VGND _1947_ net595 sg13g2_o21ai_1
XFILLER_3_306 VPWR VGND sg13g2_fill_1
XFILLER_3_339 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_28_752 VPWR VGND sg13g2_fill_1
XFILLER_27_240 VPWR VGND sg13g2_decap_4
XFILLER_16_947 VPWR VGND sg13g2_fill_1
XFILLER_43_755 VPWR VGND sg13g2_decap_8
XFILLER_24_991 VPWR VGND sg13g2_decap_8
XFILLER_3_851 VPWR VGND sg13g2_fill_2
XFILLER_2_372 VPWR VGND sg13g2_decap_8
XFILLER_3_884 VPWR VGND sg13g2_fill_1
X_2180_ _2032_ _2033_ _2034_ VPWR VGND sg13g2_nor2_1
XFILLER_19_774 VPWR VGND sg13g2_decap_8
XFILLER_19_785 VPWR VGND sg13g2_fill_1
XFILLER_30_961 VPWR VGND sg13g2_decap_8
X_3703_ _1500_ VPWR _1606_ VGND _1537_ _1605_ sg13g2_o21ai_1
X_3634_ _1538_ net780 _1539_ VPWR VGND sg13g2_nor2b_1
X_3565_ _1488_ net400 net598 VPWR VGND sg13g2_nand2_1
XFILLER_0_309 VPWR VGND sg13g2_decap_8
X_2516_ net851 _0638_ net743 _0743_ VPWR VGND _0693_ sg13g2_nand4_1
X_3496_ _1444_ net786 _0540_ VPWR VGND sg13g2_xnor2_1
X_2447_ VPWR VGND _0662_ _0673_ _0676_ net588 _0677_ _0665_ sg13g2_a221oi_1
X_2378_ _0609_ _0606_ _0608_ VPWR VGND sg13g2_nand2_1
X_4117_ net694 VGND VPWR net950 u_usb_cdc.u_ctrl_endp.state_q\[7\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_1
X_4048_ VPWR _0416_ net495 VGND sg13g2_inv_1
XFILLER_37_582 VPWR VGND sg13g2_fill_2
XFILLER_24_232 VPWR VGND sg13g2_fill_2
XFILLER_24_265 VPWR VGND sg13g2_decap_8
XFILLER_12_438 VPWR VGND sg13g2_fill_2
XFILLER_4_637 VPWR VGND sg13g2_decap_4
XFILLER_0_832 VPWR VGND sg13g2_decap_8
XFILLER_48_836 VPWR VGND sg13g2_decap_8
Xhold9 _0247_ VPWR VGND net52 sg13g2_dlygate4sd3_1
XFILLER_16_777 VPWR VGND sg13g2_decap_4
XFILLER_11_482 VPWR VGND sg13g2_fill_1
Xhold409 u_usb_cdc.u_sie.u_phy_rx.dp_q\[0\] VPWR VGND net452 sg13g2_dlygate4sd3_1
X_3350_ net816 VPWR _1346_ VGND net821 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[54\]
+ sg13g2_o21ai_1
X_2301_ _0533_ net788 VPWR VGND net785 sg13g2_nand2b_2
X_3281_ _0936_ _0937_ _1283_ VPWR VGND sg13g2_nor2b_2
XFILLER_31_4 VPWR VGND sg13g2_fill_2
X_2232_ net759 net762 _0464_ VPWR VGND sg13g2_xor2_1
X_2163_ net845 net842 net836 u_usb_cdc.u_sie.phy_state_q\[10\] _2019_ VPWR VGND sg13g2_nor4_1
XFILLER_47_880 VPWR VGND sg13g2_decap_8
XFILLER_0_1014 VPWR VGND sg13g2_decap_8
X_2094_ VPWR _1951_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[4\] VGND sg13g2_inv_1
XFILLER_34_552 VPWR VGND sg13g2_fill_2
XFILLER_34_530 VPWR VGND sg13g2_decap_8
X_2996_ _1109_ VPWR _0131_ VGND _1062_ net612 sg13g2_o21ai_1
Xclkbuf_leaf_3_clk_regs clknet_3_0__leaf_clk_regs clknet_leaf_3_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3617_ net753 _1490_ _1523_ VPWR VGND sg13g2_nor2_2
X_3548_ _0603_ _1474_ net745 _1477_ VPWR VGND sg13g2_nand3_1
XFILLER_1_629 VPWR VGND sg13g2_decap_8
X_3479_ net908 net577 _1431_ VPWR VGND sg13g2_nor2_1
XFILLER_28_46 VPWR VGND sg13g2_fill_2
XFILLER_40_544 VPWR VGND sg13g2_fill_1
XFILLER_8_217 VPWR VGND sg13g2_fill_2
XFILLER_21_791 VPWR VGND sg13g2_fill_2
XFILLER_48_633 VPWR VGND sg13g2_decap_8
XFILLER_44_872 VPWR VGND sg13g2_decap_8
X_2850_ VGND VPWR _1016_ _1020_ _1021_ _1017_ sg13g2_a21oi_1
X_2781_ net840 _0952_ _0959_ VPWR VGND sg13g2_nor2_1
Xhold217 _0245_ VPWR VGND net260 sg13g2_dlygate4sd3_1
Xhold206 _0102_ VPWR VGND net249 sg13g2_dlygate4sd3_1
X_4451_ net727 VGND VPWR net392 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[9\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_2
Xhold228 _0408_ VPWR VGND net271 sg13g2_dlygate4sd3_1
X_3402_ _1385_ _1924_ _1379_ VPWR VGND sg13g2_xnor2_1
Xhold239 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[6\] VPWR VGND net282 sg13g2_dlygate4sd3_1
X_4382_ net677 VGND VPWR _0310_ u_usb_cdc.u_sie.addr_q\[4\] clknet_leaf_50_clk_regs
+ sg13g2_dfrbpq_1
Xfanout708 _2041_ net708 VPWR VGND sg13g2_buf_8
Xfanout719 _1916_ net719 VPWR VGND sg13g2_buf_8
X_3333_ VPWR VGND _1983_ net616 _1330_ net50 _1331_ net629 sg13g2_a221oi_1
X_3264_ net829 net935 net770 _1269_ VPWR VGND sg13g2_mux2_1
X_2215_ u_usb_cdc.addr\[2\] net761 _0447_ VPWR VGND sg13g2_xor2_1
X_3195_ net342 _1222_ _1224_ VPWR VGND sg13g2_nor2_1
X_2146_ VPWR _2002_ net370 VGND sg13g2_inv_1
XFILLER_38_176 VPWR VGND sg13g2_fill_2
XFILLER_39_688 VPWR VGND sg13g2_fill_2
XFILLER_42_809 VPWR VGND sg13g2_fill_1
X_2077_ _1934_ net998 VPWR VGND sg13g2_inv_2
XFILLER_41_319 VPWR VGND sg13g2_fill_1
XFILLER_14_26 VPWR VGND sg13g2_fill_1
XFILLER_10_728 VPWR VGND sg13g2_fill_2
X_2979_ _1097_ VPWR _0123_ VGND _1040_ net612 sg13g2_o21ai_1
XFILLER_49_408 VPWR VGND sg13g2_decap_8
XFILLER_29_198 VPWR VGND sg13g2_fill_1
XFILLER_41_886 VPWR VGND sg13g2_fill_2
XFILLER_13_566 VPWR VGND sg13g2_fill_1
XFILLER_13_577 VPWR VGND sg13g2_decap_8
XFILLER_40_363 VPWR VGND sg13g2_fill_1
XFILLER_13_588 VPWR VGND sg13g2_fill_2
XFILLER_0_470 VPWR VGND sg13g2_decap_8
XFILLER_1_982 VPWR VGND sg13g2_decap_8
XFILLER_49_975 VPWR VGND sg13g2_decap_8
XFILLER_48_485 VPWR VGND sg13g2_decap_8
XFILLER_24_809 VPWR VGND sg13g2_decap_8
XFILLER_36_669 VPWR VGND sg13g2_fill_1
X_3951_ net465 net747 _1804_ VPWR VGND sg13g2_nor2_1
XFILLER_17_894 VPWR VGND sg13g2_decap_8
X_2902_ _1052_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ net645 VPWR VGND sg13g2_nand2_1
X_3882_ net361 net365 net336 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[3\] _1754_ VPWR VGND
+ sg13g2_and4_1
X_2833_ VGND VPWR net838 net594 _1006_ net261 sg13g2_a21oi_1
X_2764_ VGND VPWR _1909_ net28 _1993_ net835 sg13g2_a21oi_2
X_4503_ net702 VGND VPWR net482 _0060_ clknet_leaf_38_clk_regs sg13g2_dfrbpq_1
X_2695_ _0894_ VPWR _0895_ VGND _0650_ _0745_ sg13g2_o21ai_1
X_4434_ net731 VGND VPWR net210 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[1\] clknet_leaf_26_clk_regs
+ sg13g2_dfrbpq_1
X_4365_ net691 VGND VPWR net909 u_usb_cdc.u_ctrl_endp.max_length_q\[5\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_3316_ _1314_ VPWR _1315_ VGND net818 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[3\]
+ sg13g2_o21ai_1
X_4296_ net673 VGND VPWR net277 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[58\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_3247_ _1253_ _1983_ _1252_ VPWR VGND sg13g2_xnor2_1
X_3178_ _1215_ net146 _1213_ VPWR VGND sg13g2_nand2_1
X_2129_ VPWR _1986_ net575 VGND sg13g2_inv_1
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_42_617 VPWR VGND sg13g2_fill_2
XFILLER_41_138 VPWR VGND sg13g2_fill_1
XFILLER_10_569 VPWR VGND sg13g2_fill_1
Xhold581 u_usb_cdc.addr\[6\] VPWR VGND net900 sg13g2_dlygate4sd3_1
Xhold570 _0332_ VPWR VGND net889 sg13g2_dlygate4sd3_1
Xhold592 u_usb_cdc.u_sie.pid_q\[0\] VPWR VGND net911 sg13g2_dlygate4sd3_1
XFILLER_1_278 VPWR VGND sg13g2_fill_2
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_46_967 VPWR VGND sg13g2_decap_8
XFILLER_17_135 VPWR VGND sg13g2_fill_1
XFILLER_33_628 VPWR VGND sg13g2_fill_2
XFILLER_9_345 VPWR VGND sg13g2_decap_4
XFILLER_12_1003 VPWR VGND sg13g2_decap_8
X_2480_ _0690_ _0706_ u_usb_cdc.sie_out_data\[3\] _0708_ VPWR VGND sg13g2_nand3_1
XFILLER_49_5 VPWR VGND sg13g2_decap_8
X_4150_ net663 VGND VPWR _0079_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[4\]
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_2
X_3101_ _1167_ net111 _1151_ VPWR VGND sg13g2_nand2_1
XFILLER_1_790 VPWR VGND sg13g2_decap_8
X_4081_ _1901_ net84 _1900_ VPWR VGND sg13g2_nand2_1
XFILLER_49_772 VPWR VGND sg13g2_decap_8
X_3032_ _1124_ VPWR _0152_ VGND _1091_ _1098_ sg13g2_o21ai_1
XFILLER_37_978 VPWR VGND sg13g2_decap_8
XFILLER_36_488 VPWR VGND sg13g2_fill_1
XFILLER_24_639 VPWR VGND sg13g2_fill_2
X_3934_ _1789_ net853 _1747_ _1793_ VPWR VGND sg13g2_a21o_1
X_3865_ net496 net963 _0901_ _0368_ VPWR VGND sg13g2_mux2_1
X_2816_ _0514_ u_usb_cdc.endp\[3\] _0991_ VPWR VGND sg13g2_nor2b_1
X_3796_ _1693_ VPWR _0347_ VGND net724 net600 sg13g2_o21ai_1
X_2747_ _0932_ _0933_ _0931_ _0935_ VPWR VGND sg13g2_nand3_1
X_2678_ net710 _0511_ net841 _0880_ VPWR VGND _0522_ sg13g2_nand4_1
X_4417_ net705 VGND VPWR _0345_ u_usb_cdc.u_sie.data_q\[6\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_28_1021 VPWR VGND sg13g2_decap_8
X_4348_ net683 VGND VPWR _0276_ u_usb_cdc.u_ctrl_endp.addr_dd\[1\] clknet_leaf_49_clk_regs
+ sg13g2_dfrbpq_1
X_4279_ net658 VGND VPWR net147 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[41\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
XFILLER_28_923 VPWR VGND sg13g2_decap_8
XFILLER_43_926 VPWR VGND sg13g2_decap_8
XFILLER_35_1025 VPWR VGND sg13g2_decap_4
XFILLER_11_812 VPWR VGND sg13g2_fill_2
XFILLER_11_867 VPWR VGND sg13g2_fill_2
XFILLER_6_304 VPWR VGND sg13g2_fill_2
XFILLER_19_934 VPWR VGND sg13g2_fill_1
XFILLER_46_753 VPWR VGND sg13g2_decap_8
XFILLER_34_915 VPWR VGND sg13g2_fill_2
X_3650_ VGND VPWR net807 _1989_ _1555_ net799 sg13g2_a21oi_1
X_3581_ _0330_ net579 _0500_ net583 _1968_ VPWR VGND sg13g2_a22oi_1
X_2601_ _0820_ _0818_ _0819_ VPWR VGND sg13g2_nand2_1
X_2532_ net641 _0714_ net492 _0759_ VPWR VGND _0719_ sg13g2_nand4_1
X_2463_ _0691_ _0682_ _0689_ VPWR VGND sg13g2_nand2_1
X_4202_ net667 VGND VPWR net89 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[48\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_2394_ _0625_ u_usb_cdc.u_ctrl_endp.state_q\[7\] _0624_ VPWR VGND sg13g2_nand2_1
X_4133_ net736 VGND VPWR _0031_ u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[3\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_2
X_4064_ VGND VPWR _0923_ _1887_ _1889_ _1888_ sg13g2_a21oi_1
X_3015_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[3\]
+ net467 _1117_ _0142_ VPWR VGND sg13g2_mux2_1
XFILLER_12_609 VPWR VGND sg13g2_decap_4
XFILLER_32_491 VPWR VGND sg13g2_decap_8
XFILLER_20_642 VPWR VGND sg13g2_fill_2
X_3917_ _1780_ net437 net896 _1775_ VPWR VGND sg13g2_and3_1
XFILLER_20_664 VPWR VGND sg13g2_fill_1
X_3848_ _0899_ _1729_ net209 _1731_ VPWR VGND sg13g2_nand3_1
XFILLER_20_686 VPWR VGND sg13g2_fill_2
X_3779_ VGND VPWR net801 _1677_ _1678_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[2\]
+ sg13g2_a21oi_1
XFILLER_3_329 VPWR VGND sg13g2_fill_1
XFILLER_47_506 VPWR VGND sg13g2_decap_8
XFILLER_28_775 VPWR VGND sg13g2_fill_1
XFILLER_24_970 VPWR VGND sg13g2_decap_8
XFILLER_7_657 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_27_clk_regs clknet_3_7__leaf_clk_regs clknet_leaf_27_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_3_874 VPWR VGND sg13g2_fill_1
XFILLER_2_351 VPWR VGND sg13g2_decap_8
XFILLER_14_491 VPWR VGND sg13g2_decap_8
XFILLER_30_940 VPWR VGND sg13g2_decap_8
X_3702_ net782 VPWR _1605_ VGND net792 net785 sg13g2_o21ai_1
X_3633_ _0685_ _1537_ _1538_ VPWR VGND sg13g2_nor2_1
X_3564_ _1485_ VPWR _0321_ VGND _0867_ _1487_ sg13g2_o21ai_1
X_2515_ _0716_ _0741_ _0742_ VPWR VGND sg13g2_nor2_1
X_3495_ _1443_ net786 _1437_ VPWR VGND sg13g2_nand2_1
X_2446_ _0645_ _0675_ _0676_ VPWR VGND sg13g2_nor2_1
X_2377_ _0607_ VPWR _0608_ VGND _1928_ _0602_ sg13g2_o21ai_1
X_4116_ net694 VGND VPWR net948 u_usb_cdc.u_ctrl_endp.state_q\[6\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_29_539 VPWR VGND sg13g2_decap_8
XFILLER_17_26 VPWR VGND sg13g2_fill_2
X_4047_ _1876_ _1842_ _1875_ net642 net494 VPWR VGND sg13g2_a22oi_1
XFILLER_25_767 VPWR VGND sg13g2_decap_8
XFILLER_25_778 VPWR VGND sg13g2_fill_1
XFILLER_33_58 VPWR VGND sg13g2_decap_4
XFILLER_32_1017 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_4_616 VPWR VGND sg13g2_fill_1
XFILLER_3_115 VPWR VGND sg13g2_fill_2
XFILLER_0_811 VPWR VGND sg13g2_decap_8
XFILLER_48_815 VPWR VGND sg13g2_decap_8
XFILLER_0_888 VPWR VGND sg13g2_decap_8
XFILLER_28_561 VPWR VGND sg13g2_decap_8
XFILLER_15_233 VPWR VGND sg13g2_fill_1
XFILLER_30_214 VPWR VGND sg13g2_fill_1
XFILLER_31_737 VPWR VGND sg13g2_fill_1
XFILLER_8_922 VPWR VGND sg13g2_fill_1
XFILLER_8_999 VPWR VGND sg13g2_decap_8
X_3280_ _1264_ net826 _1282_ _0242_ VPWR VGND sg13g2_a21o_1
X_2300_ _0525_ _0526_ _0527_ _0530_ _0532_ VPWR VGND sg13g2_nor4_1
X_2231_ _0463_ u_usb_cdc.u_sie.data_q\[3\] _0462_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_815 VPWR VGND sg13g2_fill_2
XFILLER_24_4 VPWR VGND sg13g2_decap_8
X_2162_ net847 VPWR _2018_ VGND net710 _2016_ sg13g2_o21ai_1
X_2093_ VPWR _1950_ net310 VGND sg13g2_inv_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_46_391 VPWR VGND sg13g2_fill_2
XFILLER_22_715 VPWR VGND sg13g2_fill_1
X_2995_ _1109_ net88 _1108_ VPWR VGND sg13g2_nand2_1
X_3616_ _1519_ _1521_ _1518_ _1522_ VPWR VGND sg13g2_nand3_1
X_3547_ net745 VPWR _1476_ VGND _0603_ _1475_ sg13g2_o21ai_1
X_3478_ VGND VPWR net577 _1430_ _0292_ _1429_ sg13g2_a21oi_1
X_2429_ _0656_ VPWR _0659_ VGND _0542_ _0657_ sg13g2_o21ai_1
XFILLER_28_25 VPWR VGND sg13g2_decap_8
XFILLER_44_328 VPWR VGND sg13g2_fill_1
XFILLER_25_542 VPWR VGND sg13g2_decap_8
XFILLER_25_564 VPWR VGND sg13g2_fill_2
XFILLER_5_925 VPWR VGND sg13g2_decap_4
XFILLER_48_612 VPWR VGND sg13g2_decap_8
XFILLER_0_685 VPWR VGND sg13g2_decap_8
XFILLER_47_177 VPWR VGND sg13g2_fill_2
XFILLER_48_689 VPWR VGND sg13g2_decap_8
XFILLER_16_553 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_42_clk_regs clknet_3_4__leaf_clk_regs clknet_leaf_42_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2780_ net486 _0957_ _0958_ VPWR VGND sg13g2_nor2_1
XFILLER_8_763 VPWR VGND sg13g2_decap_8
Xhold207 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[16\] VPWR VGND
+ net250 sg13g2_dlygate4sd3_1
X_4450_ net727 VGND VPWR net458 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[8\] clknet_leaf_23_clk_regs
+ sg13g2_dfrbpq_1
X_4381_ net677 VGND VPWR _0309_ u_usb_cdc.u_sie.addr_q\[3\] clknet_leaf_49_clk_regs
+ sg13g2_dfrbpq_1
Xhold229 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[29\] VPWR
+ VGND net272 sg13g2_dlygate4sd3_1
Xhold218 u_usb_cdc.u_sie.addr_q\[0\] VPWR VGND net261 sg13g2_dlygate4sd3_1
X_3401_ net363 net639 u_usb_cdc.sie_in_req _1384_ VPWR VGND sg13g2_nand3_1
X_3332_ _1329_ VPWR _1330_ VGND _1288_ _1326_ sg13g2_o21ai_1
Xfanout709 _2026_ net709 VPWR VGND sg13g2_buf_8
X_3263_ _1268_ net830 _1264_ _0239_ VPWR VGND sg13g2_mux2_1
XFILLER_39_601 VPWR VGND sg13g2_decap_4
X_2214_ u_usb_cdc.addr\[1\] net762 _0446_ VPWR VGND sg13g2_xor2_1
X_3194_ VGND VPWR net723 net631 _0215_ _1223_ sg13g2_a21oi_1
XFILLER_22_1016 VPWR VGND sg13g2_decap_8
X_2145_ VPWR _2001_ net372 VGND sg13g2_inv_1
XFILLER_22_1027 VPWR VGND sg13g2_fill_2
XFILLER_39_656 VPWR VGND sg13g2_fill_2
XFILLER_38_166 VPWR VGND sg13g2_fill_1
X_2076_ VPWR _1933_ u_usb_cdc.u_sie.pid_q\[1\] VGND sg13g2_inv_1
X_2978_ VPWR _1100_ net610 VGND sg13g2_inv_1
XFILLER_22_589 VPWR VGND sg13g2_fill_2
XFILLER_2_906 VPWR VGND sg13g2_decap_8
Xhold730 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[5\] VPWR VGND net1049 sg13g2_dlygate4sd3_1
XFILLER_1_416 VPWR VGND sg13g2_decap_8
XFILLER_38_1023 VPWR VGND sg13g2_decap_4
XFILLER_13_534 VPWR VGND sg13g2_decap_4
XFILLER_13_545 VPWR VGND sg13g2_fill_2
XFILLER_40_386 VPWR VGND sg13g2_decap_8
XFILLER_45_1016 VPWR VGND sg13g2_decap_8
XFILLER_45_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_961 VPWR VGND sg13g2_decap_8
XFILLER_49_954 VPWR VGND sg13g2_decap_8
Xhold90 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[68\] VPWR VGND
+ net133 sg13g2_dlygate4sd3_1
XFILLER_48_464 VPWR VGND sg13g2_decap_8
XFILLER_35_158 VPWR VGND sg13g2_fill_1
X_3950_ _1802_ net918 _0391_ VPWR VGND sg13g2_nor2_1
XFILLER_32_821 VPWR VGND sg13g2_fill_1
X_2901_ _1051_ net119 _1037_ VPWR VGND sg13g2_nand2_1
X_3881_ _1752_ VPWR _0372_ VGND net336 _1753_ sg13g2_o21ai_1
X_2832_ _0479_ net763 _1005_ VPWR VGND net750 sg13g2_nand3b_1
X_2763_ net748 net502 _0043_ VPWR VGND sg13g2_nor2_1
X_4502_ net702 VGND VPWR _0419_ _0059_ clknet_leaf_37_clk_regs sg13g2_dfrbpq_2
X_2694_ _0894_ _0673_ _0771_ VPWR VGND sg13g2_nand2b_1
X_4433_ net735 VGND VPWR net313 u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] clknet_leaf_26_clk_regs
+ sg13g2_dfrbpq_2
X_4364_ net691 VGND VPWR _0292_ u_usb_cdc.u_ctrl_endp.max_length_q\[4\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_4295_ net675 VGND VPWR net102 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[57\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
X_3315_ VGND VPWR net818 _1996_ _1314_ net814 sg13g2_a21oi_1
XFILLER_6_1021 VPWR VGND sg13g2_decap_8
X_3246_ VGND VPWR _1981_ _1231_ _1252_ _1251_ sg13g2_a21oi_1
X_3177_ _1214_ VPWR _0207_ VGND net711 _1160_ sg13g2_o21ai_1
XFILLER_27_659 VPWR VGND sg13g2_fill_2
X_2128_ VPWR _1985_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[3\]
+ VGND sg13g2_inv_1
X_2059_ VPWR _1916_ net757 VGND sg13g2_inv_1
XFILLER_23_821 VPWR VGND sg13g2_fill_1
XFILLER_6_519 VPWR VGND sg13g2_decap_8
Xhold571 u_usb_cdc.u_sie.crc16_q\[7\] VPWR VGND net890 sg13g2_dlygate4sd3_1
Xhold560 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[7\] VPWR VGND net879 sg13g2_dlygate4sd3_1
Xhold582 u_usb_cdc.u_ctrl_endp.in_endp_q VPWR VGND net901 sg13g2_dlygate4sd3_1
Xhold593 _0355_ VPWR VGND net912 sg13g2_dlygate4sd3_1
XFILLER_18_604 VPWR VGND sg13g2_fill_1
XFILLER_46_946 VPWR VGND sg13g2_decap_8
XFILLER_18_659 VPWR VGND sg13g2_decap_8
XFILLER_45_423 VPWR VGND sg13g2_decap_8
XFILLER_25_180 VPWR VGND sg13g2_decap_4
XFILLER_40_194 VPWR VGND sg13g2_fill_1
XFILLER_5_596 VPWR VGND sg13g2_fill_2
X_3100_ _1165_ VPWR _0178_ VGND net827 _1166_ sg13g2_o21ai_1
X_4080_ _1900_ net638 _1899_ VPWR VGND sg13g2_nand2_1
XFILLER_49_751 VPWR VGND sg13g2_decap_8
XFILLER_37_902 VPWR VGND sg13g2_fill_1
XFILLER_37_913 VPWR VGND sg13g2_fill_1
X_3031_ _1124_ net139 _1118_ VPWR VGND sg13g2_nand2_1
XFILLER_32_651 VPWR VGND sg13g2_decap_4
X_3933_ net853 _1789_ _1792_ VPWR VGND sg13g2_nor2_1
X_3864_ _1739_ VPWR _1741_ VGND _2039_ net962 sg13g2_o21ai_1
XFILLER_31_161 VPWR VGND sg13g2_fill_2
X_2815_ VGND VPWR _2014_ _0990_ _0984_ _0982_ sg13g2_a21oi_2
X_3795_ net592 _1692_ net767 _1693_ VPWR VGND sg13g2_nand3_1
X_2746_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[1\] net814
+ _0934_ VPWR VGND sg13g2_xor2_1
X_2677_ VPWR _0018_ net1036 VGND sg13g2_inv_1
X_4416_ net693 VGND VPWR _0344_ u_usb_cdc.u_sie.data_q\[5\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_28_1000 VPWR VGND sg13g2_decap_8
X_4347_ net683 VGND VPWR _0275_ u_usb_cdc.u_ctrl_endp.addr_dd\[0\] clknet_leaf_49_clk_regs
+ sg13g2_dfrbpq_1
X_4278_ net658 VGND VPWR net215 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[40\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_3229_ _1242_ net129 _1156_ VPWR VGND sg13g2_nand2_1
XFILLER_43_905 VPWR VGND sg13g2_decap_8
XFILLER_28_979 VPWR VGND sg13g2_decap_8
XFILLER_35_1004 VPWR VGND sg13g2_decap_8
XFILLER_23_651 VPWR VGND sg13g2_fill_1
XFILLER_23_662 VPWR VGND sg13g2_fill_2
XFILLER_11_846 VPWR VGND sg13g2_fill_1
Xhold390 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[3\] VPWR VGND
+ net433 sg13g2_dlygate4sd3_1
XFILLER_42_1008 VPWR VGND sg13g2_decap_8
XFILLER_19_902 VPWR VGND sg13g2_fill_1
XFILLER_19_957 VPWR VGND sg13g2_decap_4
XFILLER_46_732 VPWR VGND sg13g2_decap_8
XFILLER_34_927 VPWR VGND sg13g2_fill_2
X_3580_ _0329_ net579 _0496_ _1492_ _1969_ VPWR VGND sg13g2_a22oi_1
X_2600_ u_usb_cdc.u_ctrl_endp.max_length_q\[0\] u_usb_cdc.u_ctrl_endp.max_length_q\[1\]
+ u_usb_cdc.u_ctrl_endp.max_length_q\[2\] u_usb_cdc.u_ctrl_endp.max_length_q\[3\]
+ _0819_ VPWR VGND sg13g2_nor4_1
X_2531_ _0682_ u_usb_cdc.configured_o u_usb_cdc.sie_out_data\[5\] _0758_ VPWR VGND
+ _0688_ sg13g2_nand4_1
XFILLER_6_861 VPWR VGND sg13g2_decap_8
X_2462_ _1913_ _0689_ _0690_ VPWR VGND sg13g2_and2_1
X_4201_ net678 VGND VPWR net97 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[47\]
+ clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
X_2393_ VGND VPWR u_usb_cdc.sie_in_req net640 _0624_ u_usb_cdc.sie_in_data_ack sg13g2_a21oi_1
X_4132_ net735 VGND VPWR net1008 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[2\] clknet_leaf_26_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_3_73 VPWR VGND sg13g2_fill_1
XFILLER_3_51 VPWR VGND sg13g2_fill_2
X_4063_ net835 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] _2020_ _1833_ _1888_ VPWR
+ VGND sg13g2_nor4_1
XFILLER_3_1024 VPWR VGND sg13g2_fill_1
X_3014_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net469 _1117_ _0141_ VPWR VGND sg13g2_mux2_1
X_3916_ VGND VPWR net437 _1775_ _1779_ net896 sg13g2_a21oi_1
XFILLER_20_621 VPWR VGND sg13g2_fill_2
X_3847_ _1730_ VPWR _0361_ VGND _1946_ net595 sg13g2_o21ai_1
X_3778_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[23\] u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[31\]
+ net808 _1677_ VPWR VGND sg13g2_mux2_1
X_2729_ _0922_ net308 net625 VPWR VGND sg13g2_nand2_1
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_16_905 VPWR VGND sg13g2_fill_2
XFILLER_28_798 VPWR VGND sg13g2_fill_2
XFILLER_2_330 VPWR VGND sg13g2_decap_8
XFILLER_18_1010 VPWR VGND sg13g2_decap_8
X_3701_ _1603_ VPWR _1604_ VGND _0718_ _1601_ sg13g2_o21ai_1
X_3632_ net784 _0669_ _1537_ VPWR VGND sg13g2_and2_1
XFILLER_30_996 VPWR VGND sg13g2_decap_8
XFILLER_6_680 VPWR VGND sg13g2_decap_8
X_3563_ _1487_ _0584_ _1486_ VPWR VGND sg13g2_nand2_1
X_2514_ VPWR VGND _0710_ _0738_ _0740_ _0719_ _0741_ _0731_ sg13g2_a221oi_1
X_3494_ _1437_ net789 _1442_ _0296_ VPWR VGND sg13g2_a21o_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_2445_ _0675_ net791 _1925_ VPWR VGND sg13g2_nand2_2
X_2376_ net849 net471 u_usb_cdc.u_ctrl_endp.state_q\[6\] _0607_ VPWR VGND sg13g2_nor3_1
X_4115_ net693 VGND VPWR net472 u_usb_cdc.u_ctrl_endp.state_q\[5\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
X_4046_ _1875_ _1874_ _1821_ _1834_ net459 VPWR VGND sg13g2_a22oi_1
XFILLER_25_735 VPWR VGND sg13g2_decap_8
XFILLER_37_562 VPWR VGND sg13g2_fill_2
XFILLER_37_584 VPWR VGND sg13g2_fill_1
XFILLER_40_705 VPWR VGND sg13g2_fill_2
XFILLER_20_484 VPWR VGND sg13g2_decap_4
XFILLER_21_985 VPWR VGND sg13g2_fill_2
XFILLER_0_867 VPWR VGND sg13g2_decap_8
XFILLER_16_757 VPWR VGND sg13g2_fill_1
XFILLER_23_70 VPWR VGND sg13g2_decap_4
XFILLER_11_495 VPWR VGND sg13g2_fill_2
XFILLER_8_978 VPWR VGND sg13g2_decap_8
X_2230_ _0461_ _0458_ _0462_ VPWR VGND sg13g2_xor2_1
X_2161_ net710 _2016_ _2017_ VPWR VGND sg13g2_nor2_2
X_2092_ VPWR _1949_ net209 VGND sg13g2_inv_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_34_554 VPWR VGND sg13g2_fill_1
X_2994_ _1108_ net644 _1100_ VPWR VGND sg13g2_nand2_2
XFILLER_21_226 VPWR VGND sg13g2_fill_1
XFILLER_21_237 VPWR VGND sg13g2_fill_1
XFILLER_22_749 VPWR VGND sg13g2_fill_2
XFILLER_30_771 VPWR VGND sg13g2_fill_1
X_3615_ _0761_ _1503_ net783 _1521_ VPWR VGND _1520_ sg13g2_nand4_1
X_3546_ _1475_ _1972_ _0950_ VPWR VGND sg13g2_nand2_1
X_3477_ net298 _1421_ _1430_ VPWR VGND sg13g2_nor2_1
X_2428_ net774 net781 _0658_ VPWR VGND sg13g2_nor2b_1
X_2359_ _0590_ _0565_ _0589_ VPWR VGND sg13g2_nand2b_1
XFILLER_45_808 VPWR VGND sg13g2_decap_4
X_4029_ _1860_ _1957_ net845 _1932_ net836 VPWR VGND sg13g2_a22oi_1
XFILLER_25_521 VPWR VGND sg13g2_fill_2
XFILLER_25_598 VPWR VGND sg13g2_fill_2
XFILLER_5_915 VPWR VGND sg13g2_fill_1
XFILLER_21_793 VPWR VGND sg13g2_fill_1
XFILLER_4_469 VPWR VGND sg13g2_fill_1
XFILLER_0_664 VPWR VGND sg13g2_decap_8
XFILLER_48_668 VPWR VGND sg13g2_decap_8
XFILLER_43_362 VPWR VGND sg13g2_decap_4
XFILLER_15_1024 VPWR VGND sg13g2_decap_4
Xhold208 _0099_ VPWR VGND net251 sg13g2_dlygate4sd3_1
Xhold219 _1006_ VPWR VGND net262 sg13g2_dlygate4sd3_1
X_4380_ net677 VGND VPWR net386 u_usb_cdc.u_sie.addr_q\[2\] clknet_leaf_49_clk_regs
+ sg13g2_dfrbpq_1
X_3400_ VGND VPWR _1923_ _1369_ _0261_ _1383_ sg13g2_a21oi_1
X_3331_ _1329_ _1327_ _1328_ _1324_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[2\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_4_981 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_11_clk_regs clknet_3_2__leaf_clk_regs clknet_leaf_11_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3262_ VPWR VGND _1260_ _1267_ _0714_ net755 _1268_ _1984_ sg13g2_a221oi_1
X_2213_ _0445_ net763 u_usb_cdc.addr\[0\] VPWR VGND sg13g2_xnor2_1
X_3193_ net317 net631 _1223_ VPWR VGND sg13g2_nor2_1
X_2144_ VPWR _2000_ net222 VGND sg13g2_inv_1
XFILLER_38_178 VPWR VGND sg13g2_fill_1
X_2075_ VPWR _1932_ u_usb_cdc.u_sie.pid_q\[0\] VGND sg13g2_inv_1
X_2977_ _1099_ _1041_ _1043_ VPWR VGND sg13g2_nand2_1
Xhold720 _0056_ VPWR VGND net1039 sg13g2_dlygate4sd3_1
Xhold731 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[2\] VPWR VGND net1050 sg13g2_dlygate4sd3_1
X_3529_ net381 net586 _1463_ VPWR VGND sg13g2_nor2_1
XFILLER_44_115 VPWR VGND sg13g2_fill_2
XFILLER_38_690 VPWR VGND sg13g2_fill_2
XFILLER_38_1002 VPWR VGND sg13g2_decap_8
XFILLER_26_896 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_41_888 VPWR VGND sg13g2_fill_1
XFILLER_4_255 VPWR VGND sg13g2_fill_2
XFILLER_5_789 VPWR VGND sg13g2_decap_4
XFILLER_1_940 VPWR VGND sg13g2_decap_8
XFILLER_49_933 VPWR VGND sg13g2_decap_8
XFILLER_48_443 VPWR VGND sg13g2_decap_8
Xhold80 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[67\] VPWR VGND
+ net123 sg13g2_dlygate4sd3_1
Xhold91 _0151_ VPWR VGND net134 sg13g2_dlygate4sd3_1
XFILLER_36_616 VPWR VGND sg13g2_decap_4
X_2900_ _1049_ VPWR _0094_ VGND net618 _1050_ sg13g2_o21ai_1
XFILLER_44_693 VPWR VGND sg13g2_fill_2
X_3880_ u_usb_cdc.u_sie.u_phy_rx.cnt_q\[1\] net615 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[0\]
+ _1753_ VPWR VGND sg13g2_nand3_1
X_2831_ _1004_ _1003_ net587 VPWR VGND sg13g2_nand2b_1
X_2762_ net501 _2049_ _0945_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_572 VPWR VGND sg13g2_fill_2
XFILLER_8_550 VPWR VGND sg13g2_fill_1
X_4501_ net702 VGND VPWR net309 _0058_ clknet_leaf_37_clk_regs sg13g2_dfrbpq_2
X_2693_ net573 VPWR _0029_ VGND _2043_ _0892_ sg13g2_o21ai_1
X_4432_ net699 VGND VPWR net108 u_usb_cdc.u_sie.out_eop_q clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_6_84 VPWR VGND sg13g2_fill_2
X_4363_ net691 VGND VPWR net899 u_usb_cdc.u_ctrl_endp.max_length_q\[3\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_3314_ net445 _1283_ _1313_ VPWR VGND sg13g2_nor2_1
X_4294_ net675 VGND VPWR net225 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[56\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
XFILLER_6_1000 VPWR VGND sg13g2_decap_8
X_3245_ _1251_ _1250_ _1154_ VPWR VGND sg13g2_nand2b_1
X_3176_ _1214_ net214 _1213_ VPWR VGND sg13g2_nand2_1
X_2127_ VPWR _1984_ net1003 VGND sg13g2_inv_1
X_2058_ net759 _1915_ VPWR VGND sg13g2_inv_4
XFILLER_2_726 VPWR VGND sg13g2_decap_8
Xhold561 u_usb_cdc.u_ctrl_endp.rec_q\[0\] VPWR VGND net880 sg13g2_dlygate4sd3_1
Xhold572 _0330_ VPWR VGND net891 sg13g2_dlygate4sd3_1
Xhold550 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[7\] VPWR VGND
+ net869 sg13g2_dlygate4sd3_1
Xhold594 u_usb_cdc.u_sie.crc16_q\[12\] VPWR VGND net913 sg13g2_dlygate4sd3_1
Xhold583 u_usb_cdc.u_sie.crc16_q\[3\] VPWR VGND net902 sg13g2_dlygate4sd3_1
XFILLER_46_925 VPWR VGND sg13g2_decap_8
XFILLER_18_627 VPWR VGND sg13g2_decap_8
XFILLER_18_638 VPWR VGND sg13g2_fill_1
XFILLER_14_855 VPWR VGND sg13g2_fill_2
XFILLER_14_866 VPWR VGND sg13g2_fill_1
XFILLER_41_630 VPWR VGND sg13g2_fill_1
XFILLER_49_730 VPWR VGND sg13g2_decap_8
X_3030_ _1123_ VPWR _0151_ VGND _1089_ _1098_ sg13g2_o21ai_1
X_3932_ _1791_ net717 net853 VPWR VGND sg13g2_nand2_1
X_3863_ u_usb_cdc.u_sie.u_phy_rx.rx_en_q net961 _1740_ VPWR VGND _0056_ sg13g2_nand3b_1
X_2814_ _0989_ net638 _0987_ VPWR VGND sg13g2_nand2_1
X_3794_ _1692_ _1974_ _0877_ VPWR VGND sg13g2_nand2_2
X_2745_ _0933_ net820 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[0\]
+ VPWR VGND sg13g2_xnor2_1
X_2676_ _0879_ net593 net846 net599 net837 VPWR VGND sg13g2_a22oi_1
X_4415_ net694 VGND VPWR _0343_ u_usb_cdc.u_sie.data_q\[4\] clknet_leaf_22_clk_regs
+ sg13g2_dfrbpq_2
X_4346_ net676 VGND VPWR _0274_ u_usb_cdc.addr\[6\] clknet_leaf_49_clk_regs sg13g2_dfrbpq_2
X_4277_ net657 VGND VPWR net213 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[39\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
X_3228_ _1241_ VPWR _0231_ VGND _1155_ _1178_ sg13g2_o21ai_1
XFILLER_39_251 VPWR VGND sg13g2_fill_1
X_3159_ _1205_ net257 net608 VPWR VGND sg13g2_nand2_1
XFILLER_28_958 VPWR VGND sg13g2_decap_8
XFILLER_14_107 VPWR VGND sg13g2_fill_1
XFILLER_23_685 VPWR VGND sg13g2_decap_8
XFILLER_11_869 VPWR VGND sg13g2_fill_1
XFILLER_2_523 VPWR VGND sg13g2_fill_2
Xhold380 u_usb_cdc.u_sie.u_phy_rx.stuffing_cnt_q\[1\] VPWR VGND net423 sg13g2_dlygate4sd3_1
XFILLER_2_534 VPWR VGND sg13g2_decap_8
Xhold391 _0086_ VPWR VGND net434 sg13g2_dlygate4sd3_1
XFILLER_46_711 VPWR VGND sg13g2_decap_8
XFILLER_34_917 VPWR VGND sg13g2_fill_1
XFILLER_46_788 VPWR VGND sg13g2_decap_8
XFILLER_42_994 VPWR VGND sg13g2_decap_8
XFILLER_41_482 VPWR VGND sg13g2_fill_2
X_2530_ VGND VPWR _0631_ _0756_ _0757_ _0742_ sg13g2_a21oi_1
X_2461_ _1914_ _0688_ _0689_ VPWR VGND sg13g2_and2_1
X_4200_ net668 VGND VPWR net71 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[46\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_2392_ _0623_ net743 _0617_ VPWR VGND sg13g2_nand2_1
X_4131_ net734 VGND VPWR net574 u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[1\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_3_1003 VPWR VGND sg13g2_decap_8
X_4062_ _1884_ _1886_ _1887_ VPWR VGND sg13g2_nor2_1
X_3013_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[1\]
+ net517 _1117_ _0140_ VPWR VGND sg13g2_mux2_1
XFILLER_37_777 VPWR VGND sg13g2_fill_2
XFILLER_25_939 VPWR VGND sg13g2_fill_2
X_3915_ _1777_ VPWR _0381_ VGND _1747_ _1778_ sg13g2_o21ai_1
XFILLER_20_633 VPWR VGND sg13g2_fill_2
X_3846_ _0899_ _1729_ net312 _1730_ VPWR VGND sg13g2_nand3_1
XFILLER_20_688 VPWR VGND sg13g2_fill_1
X_3777_ _1675_ VPWR _1676_ VGND net810 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[7\]
+ sg13g2_o21ai_1
X_2728_ VGND VPWR _1978_ _0918_ _0035_ _0921_ sg13g2_a21oi_1
X_2659_ _0568_ _0590_ _0868_ VPWR VGND sg13g2_nor2b_1
X_4329_ net652 VGND VPWR net1032 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[2\]
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_2
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_766 VPWR VGND sg13g2_decap_8
XFILLER_43_769 VPWR VGND sg13g2_decap_4
XFILLER_6_158 VPWR VGND sg13g2_fill_1
XFILLER_5_0 VPWR VGND sg13g2_fill_2
XFILLER_2_386 VPWR VGND sg13g2_decap_8
Xfanout690 net706 net690 VPWR VGND sg13g2_buf_8
XFILLER_19_722 VPWR VGND sg13g2_decap_8
XFILLER_19_799 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_36_clk_regs clknet_3_5__leaf_clk_regs clknet_leaf_36_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3700_ VGND VPWR u_usb_cdc.u_ctrl_endp.byte_cnt_q\[6\] _1507_ _1603_ _1602_ sg13g2_a21oi_1
XFILLER_30_975 VPWR VGND sg13g2_decap_8
X_3631_ _1536_ net560 net597 VPWR VGND sg13g2_nand2_1
X_3562_ u_usb_cdc.u_sie.in_byte_q\[0\] u_usb_cdc.u_sie.in_byte_q\[1\] net321 _1486_
+ VPWR VGND sg13g2_a21o_1
X_2513_ _0719_ _0739_ _0740_ VPWR VGND sg13g2_and2_1
XFILLER_6_692 VPWR VGND sg13g2_decap_4
X_3493_ _1439_ _1441_ _1442_ VPWR VGND sg13g2_nor2b_1
X_2444_ net788 net791 _0674_ VPWR VGND sg13g2_nor2b_1
X_2375_ net640 _0605_ _0606_ VPWR VGND sg13g2_and2_1
XFILLER_25_1004 VPWR VGND sg13g2_decap_8
X_4114_ net705 VGND VPWR _0014_ u_usb_cdc.ctrl_stall clknet_leaf_34_clk_regs sg13g2_dfrbpq_2
X_4045_ VGND VPWR _1823_ _1873_ _1874_ _1834_ sg13g2_a21oi_1
XFILLER_33_38 VPWR VGND sg13g2_fill_1
X_3829_ VPWR VGND net841 _1703_ _1715_ net1005 _1716_ _1710_ sg13g2_a221oi_1
XFILLER_21_997 VPWR VGND sg13g2_decap_8
XFILLER_3_117 VPWR VGND sg13g2_fill_1
XFILLER_3_128 VPWR VGND sg13g2_fill_1
XFILLER_47_316 VPWR VGND sg13g2_fill_2
XFILLER_28_585 VPWR VGND sg13g2_fill_2
XFILLER_8_957 VPWR VGND sg13g2_decap_8
XFILLER_48_1004 VPWR VGND sg13g2_decap_8
XFILLER_39_817 VPWR VGND sg13g2_fill_1
X_2160_ net768 u_usb_cdc.endp\[3\] u_usb_cdc.endp\[2\] _2016_ VPWR VGND sg13g2_nor3_1
X_2091_ VPWR _1948_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[3\] VGND sg13g2_inv_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_47_894 VPWR VGND sg13g2_decap_8
XFILLER_0_1028 VPWR VGND sg13g2_fill_1
XFILLER_15_780 VPWR VGND sg13g2_decap_4
XFILLER_34_599 VPWR VGND sg13g2_fill_2
X_2993_ _1107_ VPWR _0130_ VGND _1058_ net612 sg13g2_o21ai_1
X_3614_ net776 _1926_ _1520_ VPWR VGND sg13g2_nor2_2
X_3545_ net844 _0951_ _1474_ VPWR VGND sg13g2_nor2_2
X_3476_ net922 net577 _1429_ VPWR VGND sg13g2_nor2_1
X_2427_ _0657_ net780 VPWR VGND net777 sg13g2_nand2b_2
X_2358_ _0516_ _0588_ _0589_ VPWR VGND sg13g2_nor2_1
X_2289_ net753 net599 _0521_ VPWR VGND sg13g2_nor2_1
X_4028_ VGND VPWR _1859_ _1704_ _2018_ sg13g2_or2_1
XFILLER_13_728 VPWR VGND sg13g2_fill_2
XFILLER_12_238 VPWR VGND sg13g2_fill_2
XFILLER_40_558 VPWR VGND sg13g2_fill_1
XFILLER_5_949 VPWR VGND sg13g2_decap_8
XFILLER_0_643 VPWR VGND sg13g2_decap_8
XFILLER_48_647 VPWR VGND sg13g2_decap_8
XFILLER_47_179 VPWR VGND sg13g2_fill_1
XFILLER_44_886 VPWR VGND sg13g2_decap_8
XFILLER_16_588 VPWR VGND sg13g2_fill_1
Xhold209 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[1\] VPWR VGND
+ net252 sg13g2_dlygate4sd3_1
X_3330_ VGND VPWR net821 _1998_ _1328_ _1286_ sg13g2_a21oi_1
XFILLER_4_960 VPWR VGND sg13g2_decap_8
X_3261_ net755 _0601_ _1266_ _1267_ VPWR VGND sg13g2_nor3_1
Xclkbuf_leaf_51_clk_regs clknet_3_1__leaf_clk_regs clknet_leaf_51_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2212_ u_usb_cdc.addr\[3\] net760 _0444_ VPWR VGND sg13g2_xor2_1
X_3192_ net711 net826 _1175_ _1222_ VPWR VGND sg13g2_nor3_2
X_2143_ VPWR _1999_ net272 VGND sg13g2_inv_1
X_2074_ VPWR _1931_ u_usb_cdc.u_sie.out_eop_q VGND sg13g2_inv_1
XFILLER_47_691 VPWR VGND sg13g2_decap_8
XFILLER_35_875 VPWR VGND sg13g2_fill_2
X_2976_ _1098_ net740 _1041_ VPWR VGND sg13g2_nand2_2
Xhold710 _0358_ VPWR VGND net1029 sg13g2_dlygate4sd3_1
Xhold721 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_qq\[2\] VPWR VGND
+ net1040 sg13g2_dlygate4sd3_1
Xhold732 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[1\] VPWR
+ VGND net1051 sg13g2_dlygate4sd3_1
X_3528_ VGND VPWR _1915_ net585 _0310_ _1462_ sg13g2_a21oi_1
XFILLER_39_15 VPWR VGND sg13g2_fill_2
X_3459_ VGND VPWR net719 _1412_ _0287_ _1416_ sg13g2_a21oi_1
XFILLER_18_809 VPWR VGND sg13g2_fill_2
XFILLER_29_146 VPWR VGND sg13g2_fill_1
XFILLER_41_801 VPWR VGND sg13g2_decap_8
XFILLER_13_558 VPWR VGND sg13g2_fill_2
XFILLER_9_518 VPWR VGND sg13g2_decap_4
XFILLER_4_267 VPWR VGND sg13g2_fill_2
XFILLER_4_245 VPWR VGND sg13g2_fill_1
XFILLER_5_768 VPWR VGND sg13g2_fill_2
XFILLER_49_912 VPWR VGND sg13g2_decap_8
XFILLER_1_996 VPWR VGND sg13g2_decap_8
XFILLER_0_484 VPWR VGND sg13g2_decap_8
XFILLER_48_422 VPWR VGND sg13g2_decap_8
XFILLER_49_989 VPWR VGND sg13g2_decap_8
Xhold92 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[52\] VPWR VGND
+ net135 sg13g2_dlygate4sd3_1
Xhold81 _0150_ VPWR VGND net124 sg13g2_dlygate4sd3_1
Xhold70 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[37\] VPWR VGND
+ net113 sg13g2_dlygate4sd3_1
XFILLER_48_499 VPWR VGND sg13g2_decap_8
XFILLER_36_639 VPWR VGND sg13g2_decap_8
X_2830_ u_usb_cdc.addr\[0\] net594 net838 _1003_ VPWR VGND sg13g2_nand3_1
XFILLER_32_889 VPWR VGND sg13g2_fill_2
X_2761_ net748 net306 _0044_ VPWR VGND sg13g2_nor2_1
X_2692_ VGND VPWR net572 net707 _0893_ _0891_ sg13g2_a21oi_1
X_4500_ net701 VGND VPWR _0417_ _0057_ clknet_leaf_39_clk_regs sg13g2_dfrbpq_1
X_4431_ net699 VGND VPWR _0359_ u_usb_cdc.sie_out_err clknet_leaf_36_clk_regs sg13g2_dfrbpq_1
X_4362_ net691 VGND VPWR net865 u_usb_cdc.u_ctrl_endp.max_length_q\[2\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_3313_ VGND VPWR _2009_ net616 _0245_ _1312_ sg13g2_a21oi_1
XFILLER_4_790 VPWR VGND sg13g2_fill_2
X_4293_ net657 VGND VPWR _0222_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[55\]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_3244_ VGND VPWR _1250_ _1231_ _1981_ sg13g2_or2_1
X_3175_ net830 net827 net739 _1213_ VPWR VGND _1139_ sg13g2_nand4_1
X_2126_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[3\] _1983_
+ VPWR VGND sg13g2_inv_4
XFILLER_26_105 VPWR VGND sg13g2_fill_2
XFILLER_26_116 VPWR VGND sg13g2_decap_4
XFILLER_27_628 VPWR VGND sg13g2_fill_2
XFILLER_39_499 VPWR VGND sg13g2_decap_4
X_2057_ net1019 _1914_ VPWR VGND sg13g2_inv_4
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_23_834 VPWR VGND sg13g2_fill_2
X_2959_ _1086_ net198 _1079_ VPWR VGND sg13g2_nand2_1
Xhold562 u_usb_cdc.u_ctrl_endp.max_length_q\[0\] VPWR VGND net881 sg13g2_dlygate4sd3_1
Xhold551 _0090_ VPWR VGND net870 sg13g2_dlygate4sd3_1
Xhold540 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[1\] VPWR VGND
+ net859 sg13g2_dlygate4sd3_1
Xhold584 _0334_ VPWR VGND net903 sg13g2_dlygate4sd3_1
Xhold595 _0335_ VPWR VGND net914 sg13g2_dlygate4sd3_1
Xhold573 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[1\] VPWR
+ VGND net892 sg13g2_dlygate4sd3_1
XFILLER_46_904 VPWR VGND sg13g2_decap_8
XFILLER_12_1017 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_281 VPWR VGND sg13g2_decap_8
XFILLER_49_786 VPWR VGND sg13g2_decap_8
XFILLER_45_981 VPWR VGND sg13g2_decap_8
X_3931_ _1788_ VPWR _0385_ VGND _1789_ _1790_ sg13g2_o21ai_1
X_3862_ _1738_ _0889_ _0906_ _1739_ VPWR VGND sg13g2_a21o_1
X_2813_ VGND VPWR _0988_ _0978_ _0523_ sg13g2_or2_1
XFILLER_32_686 VPWR VGND sg13g2_fill_2
XFILLER_20_826 VPWR VGND sg13g2_fill_1
X_3793_ _1691_ VPWR _0346_ VGND _1689_ _1690_ sg13g2_o21ai_1
X_2744_ _0932_ net813 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[2\]
+ VPWR VGND sg13g2_xnor2_1
X_2675_ _0878_ VPWR _0028_ VGND _1974_ _0844_ sg13g2_o21ai_1
X_4414_ net693 VGND VPWR _0342_ u_usb_cdc.u_sie.data_q\[3\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_2
X_4345_ net676 VGND VPWR _0273_ u_usb_cdc.addr\[5\] clknet_leaf_48_clk_regs sg13g2_dfrbpq_2
X_4276_ net649 VGND VPWR net247 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[38\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
X_3227_ _1241_ net152 _1156_ VPWR VGND sg13g2_nand2_1
X_3158_ net711 _1153_ _1158_ _1204_ VPWR VGND sg13g2_or3_1
XFILLER_28_937 VPWR VGND sg13g2_decap_8
X_2109_ _1966_ net539 VPWR VGND sg13g2_inv_2
X_3089_ net829 _1158_ _1159_ VPWR VGND sg13g2_nor2_2
XFILLER_23_620 VPWR VGND sg13g2_fill_1
XFILLER_22_141 VPWR VGND sg13g2_decap_4
XFILLER_10_369 VPWR VGND sg13g2_fill_1
Xhold381 _1800_ VPWR VGND net424 sg13g2_dlygate4sd3_1
Xhold370 u_usb_cdc.u_ctrl_endp.dev_state_qq\[1\] VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold392 u_usb_cdc.u_ctrl_endp.addr_dd\[6\] VPWR VGND net435 sg13g2_dlygate4sd3_1
Xfanout850 u_usb_cdc.u_ctrl_endp.state_q\[2\] net850 VPWR VGND sg13g2_buf_8
XFILLER_46_767 VPWR VGND sg13g2_decap_8
XFILLER_26_60 VPWR VGND sg13g2_decap_8
XFILLER_34_929 VPWR VGND sg13g2_fill_1
XFILLER_26_491 VPWR VGND sg13g2_fill_2
XFILLER_45_288 VPWR VGND sg13g2_decap_8
XFILLER_42_973 VPWR VGND sg13g2_decap_8
XFILLER_13_130 VPWR VGND sg13g2_fill_1
XFILLER_9_101 VPWR VGND sg13g2_fill_2
X_2460_ net298 net757 u_usb_cdc.sie_out_data\[6\] _0688_ VPWR VGND sg13g2_nor3_1
XFILLER_6_874 VPWR VGND sg13g2_decap_4
X_4130_ net734 VGND VPWR net1023 _0051_ clknet_leaf_29_clk_regs sg13g2_dfrbpq_1
X_2391_ net590 _0621_ _0622_ VPWR VGND sg13g2_nor2_1
XFILLER_1_590 VPWR VGND sg13g2_decap_4
X_4061_ VGND VPWR _0059_ net308 _1886_ net481 sg13g2_a21oi_1
X_3012_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[0\]
+ net507 _1117_ _0139_ VPWR VGND sg13g2_mux2_1
XFILLER_49_583 VPWR VGND sg13g2_decap_8
XFILLER_17_491 VPWR VGND sg13g2_decap_8
X_3914_ _1778_ net437 _1775_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_984 VPWR VGND sg13g2_decap_8
X_3845_ _0912_ VPWR _1729_ VGND u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] _0905_
+ sg13g2_o21ai_1
X_3776_ VGND VPWR net810 _1992_ _1675_ net801 sg13g2_a21oi_1
X_2727_ net393 net929 _0921_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_6_clk_regs clknet_3_1__leaf_clk_regs clknet_leaf_6_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2658_ _0867_ net843 net593 VPWR VGND sg13g2_nand2_2
X_2589_ _0810_ VPWR _0010_ VGND _1942_ _0809_ sg13g2_o21ai_1
X_4328_ net652 VGND VPWR _0256_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[1\]
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
X_4259_ net654 VGND VPWR net360 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[21\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
XFILLER_43_737 VPWR VGND sg13g2_decap_4
XFILLER_42_247 VPWR VGND sg13g2_fill_1
XFILLER_24_984 VPWR VGND sg13g2_decap_8
XFILLER_7_627 VPWR VGND sg13g2_decap_8
XFILLER_12_84 VPWR VGND sg13g2_fill_2
XFILLER_2_365 VPWR VGND sg13g2_decap_8
Xfanout680 net682 net680 VPWR VGND sg13g2_buf_8
Xfanout691 net692 net691 VPWR VGND sg13g2_buf_8
XFILLER_15_940 VPWR VGND sg13g2_fill_2
XFILLER_30_954 VPWR VGND sg13g2_decap_8
X_3630_ _1497_ VPWR _0339_ VGND _1534_ _1535_ sg13g2_o21ai_1
X_3561_ _1485_ net321 net598 VPWR VGND sg13g2_nand2_1
X_2512_ _0722_ _0727_ _0739_ VPWR VGND sg13g2_nor2_1
X_3492_ _0540_ _0668_ _1441_ VPWR VGND sg13g2_nor2_2
X_2443_ net590 _0621_ net624 _0673_ VGND VPWR _0672_ sg13g2_nor4_2
X_2374_ _0605_ _0604_ _1931_ _0603_ _0602_ VPWR VGND sg13g2_a22oi_1
X_4113_ net693 VGND VPWR net970 u_usb_cdc.u_ctrl_endp.state_q\[3\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
X_4044_ _1873_ _1871_ _1872_ VPWR VGND sg13g2_nand2_1
XFILLER_37_564 VPWR VGND sg13g2_fill_1
X_3828_ VPWR _1715_ _1714_ VGND sg13g2_inv_1
XFILLER_21_987 VPWR VGND sg13g2_fill_1
X_3759_ net602 VPWR _1660_ VGND net236 _1523_ sg13g2_o21ai_1
XFILLER_0_825 VPWR VGND sg13g2_decap_8
XFILLER_48_829 VPWR VGND sg13g2_decap_8
XFILLER_16_748 VPWR VGND sg13g2_decap_4
XFILLER_43_556 VPWR VGND sg13g2_fill_1
XFILLER_23_280 VPWR VGND sg13g2_decap_4
XFILLER_24_792 VPWR VGND sg13g2_fill_1
XFILLER_7_413 VPWR VGND sg13g2_fill_2
X_2090_ VPWR _1947_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[1\] VGND sg13g2_inv_1
XFILLER_47_873 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_1007 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_34_545 VPWR VGND sg13g2_fill_2
X_2992_ _1107_ net96 _1096_ VPWR VGND sg13g2_nand2_1
XFILLER_30_762 VPWR VGND sg13g2_fill_1
X_3613_ _1519_ _1514_ u_usb_cdc.u_ctrl_endp.req_q\[2\] u_usb_cdc.configured_o u_usb_cdc.u_ctrl_endp.req_q\[4\]
+ VPWR VGND sg13g2_a22oi_1
X_3544_ net717 net1034 _1473_ _0315_ VPWR VGND sg13g2_a21o_1
X_3475_ VGND VPWR net576 _1428_ _0291_ _1427_ sg13g2_a21oi_1
X_2426_ net776 VPWR _0656_ VGND _0534_ _0655_ sg13g2_o21ai_1
XFILLER_28_39 VPWR VGND sg13g2_decap_8
X_2357_ net850 u_usb_cdc.u_ctrl_endp.state_q\[6\] _0551_ _0588_ VPWR VGND sg13g2_or3_1
X_2288_ VGND VPWR _0050_ _0519_ _0520_ net751 sg13g2_a21oi_1
X_4027_ _1858_ net292 net643 VPWR VGND sg13g2_nand2_1
XFILLER_25_523 VPWR VGND sg13g2_fill_1
XFILLER_44_38 VPWR VGND sg13g2_fill_2
XFILLER_40_526 VPWR VGND sg13g2_fill_2
XFILLER_21_784 VPWR VGND sg13g2_decap_8
XFILLER_0_611 VPWR VGND sg13g2_fill_2
XFILLER_0_622 VPWR VGND sg13g2_decap_8
XFILLER_0_699 VPWR VGND sg13g2_decap_8
XFILLER_48_626 VPWR VGND sg13g2_decap_8
XFILLER_47_114 VPWR VGND sg13g2_fill_1
XFILLER_16_512 VPWR VGND sg13g2_fill_1
XFILLER_31_526 VPWR VGND sg13g2_fill_2
XFILLER_8_733 VPWR VGND sg13g2_fill_2
X_3260_ VGND VPWR net771 _1984_ _1266_ _1265_ sg13g2_a21oi_1
X_2211_ _0443_ net758 u_usb_cdc.addr\[6\] VPWR VGND sg13g2_xnor2_1
X_3191_ _1221_ VPWR _0214_ VGND net712 _1174_ sg13g2_o21ai_1
XFILLER_22_4 VPWR VGND sg13g2_decap_8
X_2142_ VPWR _1998_ net280 VGND sg13g2_inv_1
XFILLER_38_136 VPWR VGND sg13g2_fill_2
X_2073_ VPWR _1930_ net156 VGND sg13g2_inv_1
XFILLER_35_810 VPWR VGND sg13g2_fill_1
XFILLER_47_670 VPWR VGND sg13g2_decap_8
XFILLER_35_843 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_20_clk_regs clknet_3_3__leaf_clk_regs clknet_leaf_20_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2975_ _1097_ net62 _1096_ VPWR VGND sg13g2_nand2_1
Xhold700 u_usb_cdc.sie_out_data\[5\] VPWR VGND net1019 sg13g2_dlygate4sd3_1
Xhold711 u_usb_cdc.ctrl_stall VPWR VGND net1030 sg13g2_dlygate4sd3_1
X_3527_ net408 net585 _1462_ VPWR VGND sg13g2_nor2_1
Xhold722 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[0\] VPWR
+ VGND net1041 sg13g2_dlygate4sd3_1
Xhold733 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[1\] VPWR VGND net1052 sg13g2_dlygate4sd3_1
X_3458_ net794 _1412_ _1416_ VPWR VGND sg13g2_nor2_1
XFILLER_29_103 VPWR VGND sg13g2_fill_1
X_2409_ _0639_ _0536_ _0633_ VPWR VGND sg13g2_nand2_1
X_3389_ _1374_ net809 net801 VPWR VGND sg13g2_xnor2_1
XFILLER_44_117 VPWR VGND sg13g2_fill_1
XFILLER_5_725 VPWR VGND sg13g2_decap_8
XFILLER_0_463 VPWR VGND sg13g2_decap_8
XFILLER_1_975 VPWR VGND sg13g2_decap_8
XFILLER_49_968 VPWR VGND sg13g2_decap_8
Xhold82 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[35\] VPWR VGND
+ net125 sg13g2_dlygate4sd3_1
XFILLER_29_93 VPWR VGND sg13g2_fill_1
Xhold60 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[9\] VPWR VGND
+ net103 sg13g2_dlygate4sd3_1
Xhold71 _0120_ VPWR VGND net114 sg13g2_dlygate4sd3_1
XFILLER_48_478 VPWR VGND sg13g2_decap_8
Xhold93 _0135_ VPWR VGND net136 sg13g2_dlygate4sd3_1
XFILLER_44_695 VPWR VGND sg13g2_fill_1
X_2760_ VGND VPWR u_usb_cdc.u_sie.u_phy_rx.rx_state_q\[1\] _2042_ _0944_ net305 sg13g2_a21oi_1
X_2691_ net314 VPWR _0892_ VGND _1943_ u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[3\] sg13g2_o21ai_1
XFILLER_8_574 VPWR VGND sg13g2_fill_1
X_4430_ net697 VGND VPWR net1029 u_usb_cdc.u_sie.pid_q\[3\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_6_86 VPWR VGND sg13g2_fill_1
X_4361_ net691 VGND VPWR net927 u_usb_cdc.u_ctrl_endp.max_length_q\[1\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_4292_ net673 VGND VPWR net427 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[54\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_3312_ VPWR VGND _1983_ net616 _1311_ net207 _1312_ net629 sg13g2_a221oi_1
X_3243_ net639 _0605_ net741 _1249_ VPWR VGND sg13g2_nand3_1
X_3174_ _1212_ VPWR _0206_ VGND _1192_ net609 sg13g2_o21ai_1
XFILLER_48_990 VPWR VGND sg13g2_decap_8
X_2125_ VPWR _1982_ net812 VGND sg13g2_inv_1
XFILLER_39_489 VPWR VGND sg13g2_decap_4
X_2056_ net761 _1913_ VPWR VGND sg13g2_inv_4
XFILLER_25_18 VPWR VGND sg13g2_decap_8
X_2958_ _1084_ VPWR _0117_ VGND net620 _1085_ sg13g2_o21ai_1
X_2889_ _1035_ _1042_ _1043_ VPWR VGND sg13g2_nor2_1
Xhold530 _0893_ VPWR VGND net573 sg13g2_dlygate4sd3_1
Xhold552 u_usb_cdc.u_ctrl_endp.endp_q\[1\] VPWR VGND net871 sg13g2_dlygate4sd3_1
XFILLER_9_8 VPWR VGND sg13g2_fill_1
Xhold541 _0155_ VPWR VGND net860 sg13g2_dlygate4sd3_1
Xhold563 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[3\] VPWR VGND
+ net882 sg13g2_dlygate4sd3_1
Xhold596 u_usb_cdc.u_sie.crc16_q\[8\] VPWR VGND net915 sg13g2_dlygate4sd3_1
Xhold585 u_usb_cdc.u_sie.u_phy_tx.data_q\[1\] VPWR VGND net904 sg13g2_dlygate4sd3_1
Xhold574 _0240_ VPWR VGND net893 sg13g2_dlygate4sd3_1
XFILLER_45_448 VPWR VGND sg13g2_fill_2
XFILLER_45_437 VPWR VGND sg13g2_decap_8
XFILLER_9_349 VPWR VGND sg13g2_fill_2
XFILLER_22_890 VPWR VGND sg13g2_decap_4
XFILLER_0_260 VPWR VGND sg13g2_decap_8
XFILLER_1_783 VPWR VGND sg13g2_decap_8
XFILLER_49_765 VPWR VGND sg13g2_decap_8
XFILLER_45_960 VPWR VGND sg13g2_decap_8
XFILLER_16_150 VPWR VGND sg13g2_fill_2
XFILLER_17_662 VPWR VGND sg13g2_fill_2
X_3930_ _1746_ VPWR _1790_ VGND net353 _1786_ sg13g2_o21ai_1
XFILLER_32_610 VPWR VGND sg13g2_decap_4
X_3861_ _0884_ _1737_ _0883_ _1738_ VPWR VGND sg13g2_nand3_1
X_2812_ _0523_ _0978_ _0987_ VPWR VGND sg13g2_nor2_1
X_3792_ _1691_ net984 net597 VPWR VGND sg13g2_nand2_1
X_2743_ _0931_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[3\]
+ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_q\[3\] VPWR VGND sg13g2_xnor2_1
X_2674_ _0878_ net838 net596 VPWR VGND sg13g2_nand2_1
X_4413_ net705 VGND VPWR _0341_ u_usb_cdc.u_sie.data_q\[2\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_2
X_4344_ net676 VGND VPWR _0272_ u_usb_cdc.addr\[4\] clknet_leaf_50_clk_regs sg13g2_dfrbpq_2
XFILLER_28_1014 VPWR VGND sg13g2_decap_8
X_4275_ net655 VGND VPWR net190 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[37\]
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_3226_ _1240_ VPWR _0230_ VGND net719 net604 sg13g2_o21ai_1
XFILLER_28_916 VPWR VGND sg13g2_decap_8
X_3157_ VGND VPWR _2002_ net605 _0198_ _1203_ sg13g2_a21oi_1
X_2108_ VPWR _1965_ net854 VGND sg13g2_inv_1
XFILLER_43_919 VPWR VGND sg13g2_decap_8
X_3088_ _1158_ net739 _1157_ VPWR VGND sg13g2_nand2_1
XFILLER_36_993 VPWR VGND sg13g2_decap_8
XFILLER_35_1018 VPWR VGND sg13g2_decap_8
XFILLER_23_676 VPWR VGND sg13g2_fill_2
Xhold360 _0220_ VPWR VGND net403 sg13g2_dlygate4sd3_1
Xhold371 _1471_ VPWR VGND net414 sg13g2_dlygate4sd3_1
Xhold382 _0389_ VPWR VGND net425 sg13g2_dlygate4sd3_1
Xhold393 _0281_ VPWR VGND net436 sg13g2_dlygate4sd3_1
Xfanout851 net513 net851 VPWR VGND sg13g2_buf_8
Xfanout840 net841 net840 VPWR VGND sg13g2_buf_8
XFILLER_46_746 VPWR VGND sg13g2_decap_8
XFILLER_27_982 VPWR VGND sg13g2_decap_8
XFILLER_26_83 VPWR VGND sg13g2_fill_2
XFILLER_42_952 VPWR VGND sg13g2_decap_8
XFILLER_26_94 VPWR VGND sg13g2_fill_2
XFILLER_9_113 VPWR VGND sg13g2_fill_1
XFILLER_9_179 VPWR VGND sg13g2_fill_2
XFILLER_6_886 VPWR VGND sg13g2_decap_4
X_2390_ _0609_ _0614_ _0621_ VPWR VGND _0598_ sg13g2_nand3b_1
X_4060_ _1884_ _1885_ _0419_ VPWR VGND sg13g2_nor2_1
X_3011_ VGND VPWR _1117_ net612 _1015_ sg13g2_or2_1
XFILLER_49_562 VPWR VGND sg13g2_decap_8
X_3913_ _1777_ net713 net437 VPWR VGND sg13g2_nand2_1
XFILLER_32_484 VPWR VGND sg13g2_decap_8
X_3844_ VGND VPWR _1474_ _1718_ _0360_ _1728_ sg13g2_a21oi_1
XFILLER_20_635 VPWR VGND sg13g2_fill_1
XFILLER_20_679 VPWR VGND sg13g2_decap_8
X_3775_ _1674_ VPWR _0345_ VGND _1672_ _1673_ sg13g2_o21ai_1
X_2726_ VPWR _0034_ net569 VGND sg13g2_inv_1
X_2657_ net561 VPWR _0022_ VGND _1974_ net601 sg13g2_o21ai_1
X_2588_ _0709_ _0717_ net794 _0810_ VPWR VGND _0740_ sg13g2_nand4_1
X_4327_ net648 VGND VPWR _0255_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[0\]
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_2
X_4258_ net656 VGND VPWR _0187_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[20\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_3209_ net829 net827 net831 _1231_ VPWR VGND sg13g2_nand3_1
X_4189_ net668 VGND VPWR net199 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[35\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
XFILLER_11_602 VPWR VGND sg13g2_fill_2
XFILLER_23_484 VPWR VGND sg13g2_decap_8
XFILLER_11_646 VPWR VGND sg13g2_fill_1
XFILLER_3_801 VPWR VGND sg13g2_fill_2
XFILLER_2_344 VPWR VGND sg13g2_decap_8
Xhold190 _0403_ VPWR VGND net233 sg13g2_dlygate4sd3_1
XFILLER_19_702 VPWR VGND sg13g2_decap_4
Xfanout670 net671 net670 VPWR VGND sg13g2_buf_8
Xfanout681 net682 net681 VPWR VGND sg13g2_buf_8
Xfanout692 net706 net692 VPWR VGND sg13g2_buf_8
XFILLER_19_746 VPWR VGND sg13g2_decap_4
XFILLER_37_60 VPWR VGND sg13g2_decap_8
XFILLER_15_952 VPWR VGND sg13g2_fill_2
XFILLER_30_933 VPWR VGND sg13g2_decap_8
XFILLER_18_1024 VPWR VGND sg13g2_fill_1
XFILLER_14_484 VPWR VGND sg13g2_decap_8
XFILLER_10_690 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_45_clk_regs clknet_3_4__leaf_clk_regs clknet_leaf_45_clk_regs VPWR VGND
+ sg13g2_buf_8
X_3560_ _1483_ VPWR _0320_ VGND _0867_ _1484_ sg13g2_o21ai_1
X_2511_ _0735_ _0736_ _0738_ VPWR VGND sg13g2_nor2_1
X_3491_ _1440_ VPWR _0295_ VGND net793 _1439_ sg13g2_o21ai_1
X_2442_ _0672_ _0646_ _0668_ VPWR VGND sg13g2_nand2_1
X_2373_ net755 _0601_ _0604_ VPWR VGND sg13g2_nor2_2
X_4112_ net689 VGND VPWR _0012_ u_usb_cdc.u_ctrl_endp.state_q\[2\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_2
X_4043_ VPWR VGND net842 _0570_ u_usb_cdc.u_sie.data_q\[6\] net845 _1872_ _1959_ sg13g2_a221oi_1
XFILLER_33_18 VPWR VGND sg13g2_decap_8
XFILLER_21_966 VPWR VGND sg13g2_fill_1
X_3827_ _1714_ net638 net771 net640 u_usb_cdc.ctrl_stall VPWR VGND sg13g2_a22oi_1
X_3758_ VPWR VGND _1499_ net627 _1658_ net637 _1659_ _1651_ sg13g2_a221oi_1
X_2709_ _0884_ _0907_ u_usb_cdc.u_sie.u_phy_rx.shift_register_q\[0\] _0908_ VPWR VGND
+ sg13g2_nand3_1
X_3689_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[43\] net803 _1592_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_0_804 VPWR VGND sg13g2_decap_8
XFILLER_48_808 VPWR VGND sg13g2_decap_8
XFILLER_47_318 VPWR VGND sg13g2_fill_1
XFILLER_15_226 VPWR VGND sg13g2_fill_1
XFILLER_28_587 VPWR VGND sg13g2_fill_1
XFILLER_12_966 VPWR VGND sg13g2_fill_1
XFILLER_47_852 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
X_2991_ _1106_ VPWR _0129_ VGND _1056_ net611 sg13g2_o21ai_1
XFILLER_30_741 VPWR VGND sg13g2_fill_1
X_3612_ _1512_ _1516_ _1505_ _1518_ VPWR VGND _1517_ sg13g2_nand4_1
X_3543_ net753 net717 _0436_ _0841_ _1473_ VPWR VGND sg13g2_nor4_1
X_3474_ net760 _1421_ _1428_ VPWR VGND sg13g2_nor2_1
XFILLER_43_0 VPWR VGND sg13g2_fill_2
X_2425_ _0655_ net785 net782 VPWR VGND sg13g2_nand2_1
XFILLER_28_18 VPWR VGND sg13g2_decap_8
X_2356_ _1919_ _0556_ _0564_ _0585_ _0587_ VPWR VGND sg13g2_nor4_1
X_2287_ u_usb_cdc.u_sie.phy_state_q\[2\] u_usb_cdc.u_sie.phy_state_q\[5\] u_usb_cdc.u_sie.phy_state_q\[3\]
+ _0519_ VPWR VGND sg13g2_nor3_1
X_4026_ _0413_ _1855_ _1857_ net642 _1994_ VPWR VGND sg13g2_a22oi_1
XFILLER_13_708 VPWR VGND sg13g2_fill_2
XFILLER_21_730 VPWR VGND sg13g2_fill_2
XFILLER_0_678 VPWR VGND sg13g2_decap_8
XFILLER_48_605 VPWR VGND sg13g2_decap_8
XFILLER_43_376 VPWR VGND sg13g2_fill_1
XFILLER_24_590 VPWR VGND sg13g2_decap_4
XFILLER_31_538 VPWR VGND sg13g2_fill_2
XFILLER_12_752 VPWR VGND sg13g2_fill_1
XFILLER_12_785 VPWR VGND sg13g2_fill_2
XFILLER_8_778 VPWR VGND sg13g2_decap_4
XFILLER_4_995 VPWR VGND sg13g2_decap_8
XFILLER_3_483 VPWR VGND sg13g2_fill_2
XFILLER_3_494 VPWR VGND sg13g2_fill_1
X_2210_ _0442_ net759 u_usb_cdc.addr\[4\] VPWR VGND sg13g2_xnor2_1
X_3190_ _1221_ net98 _1213_ VPWR VGND sg13g2_nand2_1
XFILLER_39_605 VPWR VGND sg13g2_fill_1
X_2141_ VPWR _1997_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[43\]
+ VGND sg13g2_inv_1
XFILLER_22_1009 VPWR VGND sg13g2_decap_8
X_2072_ _1929_ u_usb_cdc.u_ctrl_endp.state_q\[6\] VPWR VGND sg13g2_inv_2
XFILLER_35_877 VPWR VGND sg13g2_fill_1
X_2974_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\] _1985_ net740
+ _1096_ VPWR VGND net645 sg13g2_nand4_1
XFILLER_30_571 VPWR VGND sg13g2_fill_1
XFILLER_30_560 VPWR VGND sg13g2_fill_1
Xhold712 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_first_q\[2\] VPWR
+ VGND net1031 sg13g2_dlygate4sd3_1
Xhold701 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[7\]
+ VPWR VGND net1020 sg13g2_dlygate4sd3_1
X_3526_ VGND VPWR net720 net585 _0309_ _1461_ sg13g2_a21oi_1
Xhold734 u_usb_cdc.u_sie.pid_q\[2\] VPWR VGND net1053 sg13g2_dlygate4sd3_1
Xhold723 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\] VPWR
+ VGND net1042 sg13g2_dlygate4sd3_1
XFILLER_1_409 VPWR VGND sg13g2_decap_8
X_3457_ VGND VPWR _1914_ _1412_ _0286_ _1415_ sg13g2_a21oi_1
X_2408_ _0536_ _0633_ _0638_ VPWR VGND sg13g2_and2_1
X_3388_ _1373_ net811 _1369_ _0259_ VPWR VGND sg13g2_mux2_1
XFILLER_29_126 VPWR VGND sg13g2_fill_2
X_2339_ net594 _0570_ _0571_ VPWR VGND sg13g2_and2_1
X_4009_ net642 _1009_ _1842_ VPWR VGND sg13g2_nor2_2
XFILLER_26_811 VPWR VGND sg13g2_decap_8
XFILLER_38_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_1016 VPWR VGND sg13g2_decap_8
XFILLER_13_538 VPWR VGND sg13g2_fill_1
XFILLER_21_571 VPWR VGND sg13g2_decap_8
XFILLER_21_582 VPWR VGND sg13g2_fill_2
XFILLER_45_1009 VPWR VGND sg13g2_decap_8
XFILLER_1_954 VPWR VGND sg13g2_decap_8
XFILLER_0_442 VPWR VGND sg13g2_decap_8
XFILLER_48_402 VPWR VGND sg13g2_decap_8
XFILLER_49_947 VPWR VGND sg13g2_decap_8
Xhold50 _0147_ VPWR VGND net93 sg13g2_dlygate4sd3_1
Xhold83 _0202_ VPWR VGND net126 sg13g2_dlygate4sd3_1
Xhold61 _0176_ VPWR VGND net104 sg13g2_dlygate4sd3_1
Xhold72 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[15\] VPWR VGND
+ net115 sg13g2_dlygate4sd3_1
XFILLER_48_457 VPWR VGND sg13g2_decap_8
XFILLER_36_608 VPWR VGND sg13g2_fill_1
XFILLER_17_822 VPWR VGND sg13g2_fill_1
Xhold94 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[71\] VPWR VGND
+ net137 sg13g2_dlygate4sd3_1
XFILLER_12_571 VPWR VGND sg13g2_decap_8
X_2690_ VGND VPWR _2038_ _0890_ _0891_ _0881_ sg13g2_a21oi_1
X_4360_ net691 VGND VPWR _0288_ u_usb_cdc.u_ctrl_endp.max_length_q\[0\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_3311_ _1310_ VPWR _1311_ VGND _1288_ _1307_ sg13g2_o21ai_1
X_4291_ net674 VGND VPWR net403 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[53\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
XFILLER_4_792 VPWR VGND sg13g2_fill_1
X_3242_ _1248_ VPWR _0238_ VGND _1155_ _1192_ sg13g2_o21ai_1
XFILLER_39_402 VPWR VGND sg13g2_decap_8
X_3173_ _1212_ net212 net608 VPWR VGND sg13g2_nand2_1
XFILLER_6_1014 VPWR VGND sg13g2_decap_8
X_2124_ VPWR _1981_ net826 VGND sg13g2_inv_1
X_2055_ VPWR _1912_ net760 VGND sg13g2_inv_1
XFILLER_35_630 VPWR VGND sg13g2_decap_4
XFILLER_23_814 VPWR VGND sg13g2_decap_8
XFILLER_23_836 VPWR VGND sg13g2_fill_1
X_2957_ _1085_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.u_sync_data.app_in_data_q\[2\]
+ net636 VPWR VGND sg13g2_nand2_1
X_2888_ _1042_ net740 _1020_ VPWR VGND sg13g2_nand2_1
Xhold520 _0301_ VPWR VGND net563 sg13g2_dlygate4sd3_1
Xhold531 _0029_ VPWR VGND net574 sg13g2_dlygate4sd3_1
Xhold542 u_usb_cdc.addr\[2\] VPWR VGND net861 sg13g2_dlygate4sd3_1
Xhold553 u_usb_cdc.u_sie.u_phy_tx.tx_state_q\[2\] VPWR VGND net872 sg13g2_dlygate4sd3_1
Xhold575 u_usb_cdc.u_ctrl_endp.req_q\[1\] VPWR VGND net894 sg13g2_dlygate4sd3_1
Xhold586 u_usb_cdc.addr\[1\] VPWR VGND net905 sg13g2_dlygate4sd3_1
Xhold597 _0331_ VPWR VGND net916 sg13g2_dlygate4sd3_1
X_4489_ net733 VGND VPWR net13 u_usb_cdc.u_sie.u_phy_rx.dp_q\[2\] clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_1
Xhold564 _0157_ VPWR VGND net883 sg13g2_dlygate4sd3_1
X_3509_ _1449_ net774 _1454_ VPWR VGND sg13g2_xor2_1
XFILLER_46_939 VPWR VGND sg13g2_decap_8
XFILLER_26_641 VPWR VGND sg13g2_fill_2
XFILLER_25_173 VPWR VGND sg13g2_decap_8
XFILLER_25_184 VPWR VGND sg13g2_fill_2
XFILLER_9_317 VPWR VGND sg13g2_fill_1
XFILLER_5_501 VPWR VGND sg13g2_fill_1
XFILLER_5_523 VPWR VGND sg13g2_fill_2
XFILLER_1_762 VPWR VGND sg13g2_decap_8
XFILLER_49_744 VPWR VGND sg13g2_decap_8
XFILLER_44_460 VPWR VGND sg13g2_fill_2
X_3860_ _1737_ _0056_ _1946_ VPWR VGND sg13g2_nand2_1
XFILLER_32_644 VPWR VGND sg13g2_decap_8
X_2811_ _0981_ VPWR _0069_ VGND _0980_ _0986_ sg13g2_o21ai_1
X_3791_ _0439_ VPWR _1690_ VGND net270 _1523_ sg13g2_o21ai_1
X_2742_ net61 net49 _0041_ VPWR VGND sg13g2_and2_1
XFILLER_9_884 VPWR VGND sg13g2_fill_2
X_2673_ _0876_ VPWR _0027_ VGND _0844_ _0877_ sg13g2_o21ai_1
X_4412_ net706 VGND VPWR _0340_ u_usb_cdc.u_sie.data_q\[1\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_2
X_4343_ net683 VGND VPWR _0271_ u_usb_cdc.addr\[3\] clknet_leaf_49_clk_regs sg13g2_dfrbpq_2
X_4274_ net654 VGND VPWR net186 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[36\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_3225_ _1240_ net148 net604 VPWR VGND sg13g2_nand2_1
X_3156_ net757 net606 _1203_ VPWR VGND sg13g2_nor2_1
X_3087_ _1157_ net826 _1154_ VPWR VGND sg13g2_xnor2_1
X_2107_ VPWR _1964_ net902 VGND sg13g2_inv_1
XFILLER_23_611 VPWR VGND sg13g2_decap_8
XFILLER_10_305 VPWR VGND sg13g2_fill_1
X_3989_ _1824_ net767 net842 u_usb_cdc.u_sie.pid_q\[0\] u_usb_cdc.u_sie.phy_state_q\[11\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_22_198 VPWR VGND sg13g2_fill_2
XFILLER_2_548 VPWR VGND sg13g2_fill_2
Xhold361 u_usb_cdc.u_sie.u_phy_tx.stuffing_cnt_q\[2\] VPWR VGND net404 sg13g2_dlygate4sd3_1
Xhold350 u_usb_cdc.u_sie.u_phy_rx.state_q\[1\] VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold383 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[54\] VPWR
+ VGND net426 sg13g2_dlygate4sd3_1
Xhold372 _0314_ VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold394 u_usb_cdc.u_sie.u_phy_rx.cnt_q\[11\] VPWR VGND net437 sg13g2_dlygate4sd3_1
Xfanout841 net1017 net841 VPWR VGND sg13g2_buf_8
Xfanout830 net832 net830 VPWR VGND sg13g2_buf_8
Xdelaybuf_0_clk delaynet_0_clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_46_725 VPWR VGND sg13g2_decap_8
XFILLER_27_961 VPWR VGND sg13g2_decap_8
XFILLER_42_931 VPWR VGND sg13g2_decap_8
XFILLER_26_493 VPWR VGND sg13g2_fill_1
XFILLER_9_103 VPWR VGND sg13g2_fill_1
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_22 VPWR VGND sg13g2_fill_2
XFILLER_49_541 VPWR VGND sg13g2_decap_8
XFILLER_3_1017 VPWR VGND sg13g2_decap_8
X_3010_ _1116_ VPWR _0138_ VGND _1076_ net612 sg13g2_o21ai_1
XFILLER_36_257 VPWR VGND sg13g2_fill_2
XFILLER_45_780 VPWR VGND sg13g2_decap_8
X_3912_ _1774_ VPWR _0380_ VGND _1775_ _1776_ sg13g2_o21ai_1
X_3843_ VGND VPWR _1725_ _1727_ _1728_ net107 sg13g2_a21oi_1
X_3774_ _1674_ net992 net597 VPWR VGND sg13g2_nand2_1
X_2725_ _0920_ _0917_ net568 _2006_ net744 VPWR VGND sg13g2_a22oi_1
X_2656_ net766 _0845_ _0863_ _0866_ VPWR VGND sg13g2_or3_1
X_2587_ VGND VPWR _0641_ net622 _0809_ _0678_ sg13g2_a21oi_1
X_4326_ net652 VGND VPWR net544 u_usb_cdc.out_valid_o[0] clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
XFILLER_41_1012 VPWR VGND sg13g2_decap_8
X_4257_ net656 VGND VPWR net332 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[19\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
XFILLER_47_28 VPWR VGND sg13g2_decap_8
X_3208_ VGND VPWR net719 net631 _0222_ _1230_ sg13g2_a21oi_1
X_4188_ net666 VGND VPWR net155 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[34\]
+ clknet_leaf_7_clk_regs sg13g2_dfrbpq_1
X_3139_ _1193_ net830 net829 VPWR VGND sg13g2_nand2_2
XFILLER_24_920 VPWR VGND sg13g2_fill_1
XFILLER_6_117 VPWR VGND sg13g2_fill_2
Xhold180 _0181_ VPWR VGND net223 sg13g2_dlygate4sd3_1
XFILLER_3_868 VPWR VGND sg13g2_fill_2
Xhold191 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[46\] VPWR
+ VGND net234 sg13g2_dlygate4sd3_1
Xfanout660 net661 net660 VPWR VGND sg13g2_buf_8
Xfanout693 net694 net693 VPWR VGND sg13g2_buf_8
Xfanout671 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.rstn net671 VPWR VGND sg13g2_buf_8
Xfanout682 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.rstn net682 VPWR VGND sg13g2_buf_8
XFILLER_19_736 VPWR VGND sg13g2_decap_4
XFILLER_30_912 VPWR VGND sg13g2_decap_8
XFILLER_30_989 VPWR VGND sg13g2_decap_8
Xclkbuf_3_7__f_clk_regs clknet_0_clk_regs clknet_3_7__leaf_clk_regs VPWR VGND sg13g2_buf_8
X_2510_ VPWR _0737_ _0736_ VGND sg13g2_inv_1
X_3490_ _1440_ net793 _1437_ VPWR VGND sg13g2_nand2_1
X_2441_ _0645_ _0669_ _0671_ VPWR VGND sg13g2_nor2_1
X_2372_ net430 net354 net156 _0603_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_14_clk_regs clknet_3_2__leaf_clk_regs clknet_leaf_14_clk_regs VPWR VGND
+ sg13g2_buf_8
X_4111_ net693 VGND VPWR net960 u_usb_cdc.u_ctrl_endp.state_q\[1\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_25_1018 VPWR VGND sg13g2_decap_8
X_4042_ _1871_ _1963_ net837 _1934_ net836 VPWR VGND sg13g2_a22oi_1
XFILLER_49_360 VPWR VGND sg13g2_decap_8
X_3826_ _1713_ net848 _1712_ VPWR VGND sg13g2_nand2b_1
XFILLER_20_488 VPWR VGND sg13g2_fill_2
X_3757_ _1653_ VPWR _1658_ VGND _1655_ _1657_ sg13g2_o21ai_1
X_2708_ VGND VPWR _2037_ _0882_ _0907_ _0906_ sg13g2_a21oi_1
X_3688_ _1590_ VPWR _1591_ VGND net799 _1588_ sg13g2_o21ai_1
X_2639_ u_usb_cdc.u_sie.addr_q\[0\] u_usb_cdc.addr\[0\] _0850_ VPWR VGND sg13g2_xor2_1
X_4309_ net650 VGND VPWR net171 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[71\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
XFILLER_28_599 VPWR VGND sg13g2_decap_8
XFILLER_8_905 VPWR VGND sg13g2_fill_2
XFILLER_24_783 VPWR VGND sg13g2_decap_4
XFILLER_7_415 VPWR VGND sg13g2_fill_1
XFILLER_48_1018 VPWR VGND sg13g2_decap_8
XFILLER_47_831 VPWR VGND sg13g2_decap_8
XFILLER_19_544 VPWR VGND sg13g2_fill_2
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_19_599 VPWR VGND sg13g2_fill_1
XFILLER_34_547 VPWR VGND sg13g2_fill_1
XFILLER_15_761 VPWR VGND sg13g2_fill_2
X_2990_ _1106_ net70 _1096_ VPWR VGND sg13g2_nand2_1
XFILLER_14_282 VPWR VGND sg13g2_fill_2
X_3611_ VGND VPWR _1510_ _1511_ _1517_ _1509_ sg13g2_a21oi_1
XFILLER_30_786 VPWR VGND sg13g2_fill_1
X_3542_ net414 VPWR _0314_ VGND _1466_ _1472_ sg13g2_o21ai_1
XFILLER_7_993 VPWR VGND sg13g2_decap_8
X_3473_ net898 net576 _1427_ VPWR VGND sg13g2_nor2_1
X_2424_ net777 _0653_ _0654_ VPWR VGND sg13g2_nor2_1
XFILLER_9_1023 VPWR VGND sg13g2_decap_4
X_2355_ _1919_ _0585_ _0586_ VPWR VGND sg13g2_nor2_1
XFILLER_38_820 VPWR VGND sg13g2_fill_1
X_2286_ u_usb_cdc.ctrl_stall net640 net847 _0518_ VPWR VGND sg13g2_nand3_1
XFILLER_38_875 VPWR VGND sg13g2_fill_1
X_4025_ VGND VPWR net292 _1856_ _1857_ net642 sg13g2_a21oi_1
X_3809_ net592 _1692_ net984 _1700_ VPWR VGND sg13g2_nand3_1
XFILLER_0_657 VPWR VGND sg13g2_decap_8
XFILLER_43_333 VPWR VGND sg13g2_fill_1
XFILLER_43_366 VPWR VGND sg13g2_fill_1
XFILLER_31_528 VPWR VGND sg13g2_fill_1
XFILLER_12_764 VPWR VGND sg13g2_decap_4
XFILLER_15_1017 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_285 VPWR VGND sg13g2_fill_1
XFILLER_4_974 VPWR VGND sg13g2_decap_8
X_2140_ VPWR _1996_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[11\]
+ VGND sg13g2_inv_1
XFILLER_38_116 VPWR VGND sg13g2_fill_2
X_2071_ VPWR _1928_ net949 VGND sg13g2_inv_1
XFILLER_38_138 VPWR VGND sg13g2_fill_1
XFILLER_22_539 VPWR VGND sg13g2_decap_4
X_2973_ _1094_ VPWR _0122_ VGND net620 _1095_ sg13g2_o21ai_1
Xhold702 u_usb_cdc.u_ctrl_endp.byte_cnt_q\[4\] VPWR VGND net1021 sg13g2_dlygate4sd3_1
X_3525_ net448 net585 _1461_ VPWR VGND sg13g2_nor2_1
Xhold735 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_last_qq\[3\] VPWR
+ VGND net1054 sg13g2_dlygate4sd3_1
Xhold713 _0257_ VPWR VGND net1032 sg13g2_dlygate4sd3_1
Xhold724 u_usb_cdc.sie_out_err VPWR VGND net1043 sg13g2_dlygate4sd3_1
X_3456_ net492 _1412_ _1415_ VPWR VGND sg13g2_nor2_1
X_2407_ _0611_ _0616_ net624 _0637_ VGND VPWR _0636_ sg13g2_nor4_2
X_3387_ _1370_ VPWR _1373_ VGND net809 _1372_ sg13g2_o21ai_1
X_2338_ _2017_ _0569_ _0570_ VPWR VGND sg13g2_nor2_1
X_2269_ _0501_ net915 u_usb_cdc.u_sie.data_q\[7\] VPWR VGND sg13g2_xnor2_1
X_4008_ net642 net904 _1841_ _0411_ VPWR VGND sg13g2_a21o_1
XFILLER_26_889 VPWR VGND sg13g2_decap_8
XFILLER_0_421 VPWR VGND sg13g2_decap_8
XFILLER_1_933 VPWR VGND sg13g2_decap_8
XFILLER_49_926 VPWR VGND sg13g2_decap_8
XFILLER_0_498 VPWR VGND sg13g2_decap_8
Xhold40 _0091_ VPWR VGND net83 sg13g2_dlygate4sd3_1
XFILLER_48_436 VPWR VGND sg13g2_decap_8
Xhold73 _0182_ VPWR VGND net116 sg13g2_dlygate4sd3_1
Xhold51 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[20\] VPWR VGND
+ net94 sg13g2_dlygate4sd3_1
Xhold62 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_fifo_q\[15\] VPWR VGND
+ net105 sg13g2_dlygate4sd3_1
Xhold84 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[43\] VPWR VGND
+ net127 sg13g2_dlygate4sd3_1
XFILLER_29_683 VPWR VGND sg13g2_fill_1
XFILLER_35_108 VPWR VGND sg13g2_fill_2
Xhold95 _0154_ VPWR VGND net138 sg13g2_dlygate4sd3_1
XFILLER_28_171 VPWR VGND sg13g2_fill_2
XFILLER_17_878 VPWR VGND sg13g2_fill_2
XFILLER_44_686 VPWR VGND sg13g2_decap_8
X_3310_ _1310_ _1308_ _1309_ _1305_ net812 VPWR VGND sg13g2_a22oi_1
X_4290_ net672 VGND VPWR _0219_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[52\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
XFILLER_3_292 VPWR VGND sg13g2_fill_2
X_3241_ _1248_ net170 _1156_ VPWR VGND sg13g2_nand2_1
X_3172_ _1211_ VPWR _0205_ VGND _1190_ net609 sg13g2_o21ai_1
X_2123_ VPWR _1980_ net828 VGND sg13g2_inv_1
XFILLER_39_447 VPWR VGND sg13g2_fill_2
X_2054_ VPWR _1911_ net762 VGND sg13g2_inv_1
XFILLER_23_804 VPWR VGND sg13g2_fill_1
XFILLER_35_675 VPWR VGND sg13g2_decap_4
X_2956_ _1084_ net154 _1079_ VPWR VGND sg13g2_nand2_1
X_2887_ _1018_ u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_q\[2\] _1041_
+ VPWR VGND sg13g2_xor2_1
Xhold510 u_usb_cdc.u_sie.u_phy_rx.nrzi_q\[0\] VPWR VGND net553 sg13g2_dlygate4sd3_1
XFILLER_2_719 VPWR VGND sg13g2_decap_8
Xhold521 u_usb_cdc.u_ctrl_endp.max_length_q\[6\] VPWR VGND net564 sg13g2_dlygate4sd3_1
Xhold554 _2029_ VPWR VGND net873 sg13g2_dlygate4sd3_1
Xhold543 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[2\] VPWR VGND
+ net862 sg13g2_dlygate4sd3_1
Xhold532 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_first_q\[1\] VPWR VGND
+ net575 sg13g2_dlygate4sd3_1
Xhold576 _0002_ VPWR VGND net895 sg13g2_dlygate4sd3_1
Xhold587 u_usb_cdc.u_sie.crc16_q\[6\] VPWR VGND net906 sg13g2_dlygate4sd3_1
X_4488_ net733 VGND VPWR net46 u_usb_cdc.u_sie.u_phy_rx.dp_q\[1\] clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_1
Xhold565 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_in_fifo.in_last_qq\[0\] VPWR VGND
+ net884 sg13g2_dlygate4sd3_1
X_3508_ _1446_ _1452_ _1453_ VPWR VGND sg13g2_nor2_1
X_3439_ VGND VPWR net720 net582 _0278_ _1405_ sg13g2_a21oi_1
Xhold598 u_usb_cdc.bus_reset VPWR VGND net917 sg13g2_dlygate4sd3_1
XFILLER_46_918 VPWR VGND sg13g2_decap_8
XFILLER_39_981 VPWR VGND sg13g2_decap_8
XFILLER_38_491 VPWR VGND sg13g2_decap_8
XFILLER_25_130 VPWR VGND sg13g2_decap_8
XFILLER_25_152 VPWR VGND sg13g2_decap_8
Xoutput30 net30 usb_dp_tx_o VPWR VGND sg13g2_buf_1
XFILLER_1_741 VPWR VGND sg13g2_decap_8
XFILLER_49_723 VPWR VGND sg13g2_decap_8
XFILLER_0_295 VPWR VGND sg13g2_decap_8
XFILLER_17_631 VPWR VGND sg13g2_fill_1
XFILLER_45_995 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_39_clk_regs clknet_3_5__leaf_clk_regs clknet_leaf_39_clk_regs VPWR VGND
+ sg13g2_buf_8
X_2810_ net838 _0985_ _0986_ VPWR VGND sg13g2_nor2_1
X_3790_ VPWR VGND _1499_ net627 _1688_ net637 _1689_ _1686_ sg13g2_a221oi_1
XFILLER_32_678 VPWR VGND sg13g2_fill_2
X_2741_ _0929_ VPWR _0003_ VGND _0632_ _0930_ sg13g2_o21ai_1
XFILLER_8_373 VPWR VGND sg13g2_fill_1
XFILLER_8_340 VPWR VGND sg13g2_decap_8
X_2672_ net841 net524 _0877_ VPWR VGND sg13g2_nor2_2
X_4411_ net705 VGND VPWR _0339_ u_usb_cdc.u_sie.data_q\[0\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_2
X_4342_ net676 VGND VPWR _0270_ u_usb_cdc.addr\[2\] clknet_leaf_47_clk_regs sg13g2_dfrbpq_2
X_4273_ net649 VGND VPWR net126 u_usb_cdc.u_bulk_endps\[0\].u_bulk_endp.u_out_fifo.out_fifo_q\[35\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
X_3224_ VGND VPWR _2001_ net603 _0229_ _1239_ sg13g2_a21oi_1
.ends

