magic
tech ihp-sg13g2
magscale 1 2
timestamp 1755175755
<< metal1 >>
rect 576 13628 14400 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 14400 13628
rect 576 13564 14400 13588
rect 5259 13376 5301 13385
rect 5259 13336 5260 13376
rect 5300 13336 5301 13376
rect 5259 13327 5301 13336
rect 6891 13376 6933 13385
rect 6891 13336 6892 13376
rect 6932 13336 6933 13376
rect 6891 13327 6933 13336
rect 11211 13376 11253 13385
rect 11211 13336 11212 13376
rect 11252 13336 11253 13376
rect 11211 13327 11253 13336
rect 7075 13208 7133 13209
rect 7075 13168 7084 13208
rect 7124 13168 7133 13208
rect 7075 13167 7133 13168
rect 7179 13208 7221 13217
rect 7179 13168 7180 13208
rect 7220 13168 7221 13208
rect 7179 13159 7221 13168
rect 7371 13208 7413 13217
rect 7371 13168 7372 13208
rect 7412 13168 7413 13208
rect 7371 13159 7413 13168
rect 8227 13208 8285 13209
rect 8227 13168 8236 13208
rect 8276 13168 8285 13208
rect 8227 13167 8285 13168
rect 8811 13208 8853 13217
rect 8811 13168 8812 13208
rect 8852 13168 8853 13208
rect 8811 13159 8853 13168
rect 8907 13208 8949 13217
rect 8907 13168 8908 13208
rect 8948 13168 8949 13208
rect 8907 13159 8949 13168
rect 9483 13208 9525 13217
rect 9483 13168 9484 13208
rect 9524 13168 9525 13208
rect 9483 13159 9525 13168
rect 10147 13208 10205 13209
rect 10147 13168 10156 13208
rect 10196 13168 10205 13208
rect 10147 13167 10205 13168
rect 10347 13208 10389 13217
rect 10347 13168 10348 13208
rect 10388 13168 10389 13208
rect 10347 13159 10389 13168
rect 10539 13208 10581 13217
rect 10539 13168 10540 13208
rect 10580 13168 10581 13208
rect 10539 13159 10581 13168
rect 10915 13208 10973 13209
rect 10915 13168 10924 13208
rect 10964 13168 10973 13208
rect 10915 13167 10973 13168
rect 12355 13208 12413 13209
rect 12355 13168 12364 13208
rect 12404 13168 12413 13208
rect 12355 13167 12413 13168
rect 9091 13124 9149 13125
rect 9091 13084 9100 13124
rect 9140 13084 9149 13124
rect 9091 13083 9149 13084
rect 7267 13040 7325 13041
rect 7267 13000 7276 13040
rect 7316 13000 7325 13040
rect 7267 12999 7325 13000
rect 7555 13040 7613 13041
rect 7555 13000 7564 13040
rect 7604 13000 7613 13040
rect 7555 12999 7613 13000
rect 8803 13040 8861 13041
rect 8803 13000 8812 13040
rect 8852 13000 8861 13040
rect 8803 12999 8861 13000
rect 10443 13040 10485 13049
rect 10443 13000 10444 13040
rect 10484 13000 10485 13040
rect 10443 12991 10485 13000
rect 10723 13040 10781 13041
rect 10723 13000 10732 13040
rect 10772 13000 10781 13040
rect 10723 12999 10781 13000
rect 11011 13040 11069 13041
rect 11011 13000 11020 13040
rect 11060 13000 11069 13040
rect 11011 12999 11069 13000
rect 11683 13040 11741 13041
rect 11683 13000 11692 13040
rect 11732 13000 11741 13040
rect 11683 12999 11741 13000
rect 576 12872 14400 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 14400 12872
rect 576 12808 14400 12832
rect 7659 12704 7701 12713
rect 7659 12664 7660 12704
rect 7700 12664 7701 12704
rect 7659 12655 7701 12664
rect 8427 12620 8469 12629
rect 8427 12580 8428 12620
rect 8468 12580 8469 12620
rect 8427 12571 8469 12580
rect 3427 12536 3485 12537
rect 3427 12496 3436 12536
rect 3476 12496 3485 12536
rect 3427 12495 3485 12496
rect 4771 12536 4829 12537
rect 4771 12496 4780 12536
rect 4820 12496 4829 12536
rect 4771 12495 4829 12496
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 4971 12487 5013 12496
rect 5259 12536 5301 12545
rect 5259 12496 5260 12536
rect 5300 12496 5301 12536
rect 5259 12487 5301 12496
rect 5451 12536 5493 12545
rect 5451 12496 5452 12536
rect 5492 12496 5493 12536
rect 5451 12487 5493 12496
rect 6115 12536 6173 12537
rect 6115 12496 6124 12536
rect 6164 12496 6173 12536
rect 6115 12495 6173 12496
rect 7275 12536 7317 12545
rect 7275 12496 7276 12536
rect 7316 12496 7317 12536
rect 7275 12487 7317 12496
rect 7467 12536 7509 12545
rect 7467 12496 7468 12536
rect 7508 12496 7509 12536
rect 7467 12487 7509 12496
rect 7843 12536 7901 12537
rect 7843 12496 7852 12536
rect 7892 12496 7901 12536
rect 7843 12495 7901 12496
rect 7939 12536 7997 12537
rect 7939 12496 7948 12536
rect 7988 12496 7997 12536
rect 7939 12495 7997 12496
rect 9091 12536 9149 12537
rect 9091 12496 9100 12536
rect 9140 12496 9149 12536
rect 9091 12495 9149 12496
rect 9955 12536 10013 12537
rect 9955 12496 9964 12536
rect 10004 12496 10013 12536
rect 9955 12495 10013 12496
rect 10347 12536 10389 12545
rect 10347 12496 10348 12536
rect 10388 12496 10389 12536
rect 10347 12487 10389 12496
rect 10723 12536 10781 12537
rect 10723 12496 10732 12536
rect 10772 12496 10781 12536
rect 10723 12495 10781 12496
rect 11587 12536 11645 12537
rect 11587 12496 11596 12536
rect 11636 12496 11645 12536
rect 11587 12495 11645 12496
rect 1131 12368 1173 12377
rect 1131 12328 1132 12368
rect 1172 12328 1173 12368
rect 1131 12319 1173 12328
rect 2571 12368 2613 12377
rect 2571 12328 2572 12368
rect 2612 12328 2613 12368
rect 2571 12319 2613 12328
rect 3723 12368 3765 12377
rect 3723 12328 3724 12368
rect 3764 12328 3765 12368
rect 3723 12319 3765 12328
rect 6795 12368 6837 12377
rect 6795 12328 6796 12368
rect 6836 12328 6837 12368
rect 6795 12319 6837 12328
rect 12939 12368 12981 12377
rect 12939 12328 12940 12368
rect 12980 12328 12981 12368
rect 12939 12319 12981 12328
rect 2755 12284 2813 12285
rect 2755 12244 2764 12284
rect 2804 12244 2813 12284
rect 2755 12243 2813 12244
rect 4099 12284 4157 12285
rect 4099 12244 4108 12284
rect 4148 12244 4157 12284
rect 4099 12243 4157 12244
rect 5259 12284 5301 12293
rect 5259 12244 5260 12284
rect 5300 12244 5301 12284
rect 5259 12235 5301 12244
rect 7275 12284 7317 12293
rect 7275 12244 7276 12284
rect 7316 12244 7317 12284
rect 7275 12235 7317 12244
rect 9283 12284 9341 12285
rect 9283 12244 9292 12284
rect 9332 12244 9341 12284
rect 9283 12243 9341 12244
rect 12739 12284 12797 12285
rect 12739 12244 12748 12284
rect 12788 12244 12797 12284
rect 12739 12243 12797 12244
rect 576 12116 14400 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 14400 12116
rect 576 12052 14400 12076
rect 3043 11948 3101 11949
rect 3043 11908 3052 11948
rect 3092 11908 3101 11948
rect 3043 11907 3101 11908
rect 5731 11948 5789 11949
rect 5731 11908 5740 11948
rect 5780 11908 5789 11948
rect 5731 11907 5789 11908
rect 8715 11864 8757 11873
rect 8715 11824 8716 11864
rect 8756 11824 8757 11864
rect 8715 11815 8757 11824
rect 1027 11696 1085 11697
rect 1027 11656 1036 11696
rect 1076 11656 1085 11696
rect 1027 11655 1085 11656
rect 1891 11696 1949 11697
rect 1891 11656 1900 11696
rect 1940 11656 1949 11696
rect 1891 11655 1949 11656
rect 3339 11696 3381 11705
rect 3339 11656 3340 11696
rect 3380 11656 3381 11696
rect 3339 11647 3381 11656
rect 3715 11696 3773 11697
rect 3715 11656 3724 11696
rect 3764 11656 3773 11696
rect 3715 11655 3773 11656
rect 4579 11696 4637 11697
rect 4579 11656 4588 11696
rect 4628 11656 4637 11696
rect 4579 11655 4637 11656
rect 6315 11696 6357 11705
rect 6315 11656 6316 11696
rect 6356 11656 6357 11696
rect 6315 11647 6357 11656
rect 6691 11696 6749 11697
rect 6691 11656 6700 11696
rect 6740 11656 6749 11696
rect 6691 11655 6749 11656
rect 7555 11696 7613 11697
rect 7555 11656 7564 11696
rect 7604 11656 7613 11696
rect 7555 11655 7613 11656
rect 9667 11696 9725 11697
rect 9667 11656 9676 11696
rect 9716 11656 9725 11696
rect 9667 11655 9725 11656
rect 10059 11696 10101 11705
rect 10059 11656 10060 11696
rect 10100 11656 10101 11696
rect 10059 11647 10101 11656
rect 10147 11696 10205 11697
rect 10147 11656 10156 11696
rect 10196 11656 10205 11696
rect 10147 11655 10205 11656
rect 10827 11696 10869 11705
rect 10827 11656 10828 11696
rect 10868 11656 10869 11696
rect 10827 11647 10869 11656
rect 11683 11696 11741 11697
rect 11683 11656 11692 11696
rect 11732 11656 11741 11696
rect 11683 11655 11741 11656
rect 12259 11696 12317 11697
rect 12259 11656 12268 11696
rect 12308 11656 12317 11696
rect 12259 11655 12317 11656
rect 13123 11696 13181 11697
rect 13123 11656 13132 11696
rect 13172 11656 13181 11696
rect 13123 11655 13181 11656
rect 651 11612 693 11621
rect 651 11572 652 11612
rect 692 11572 693 11612
rect 651 11563 693 11572
rect 11883 11612 11925 11621
rect 11883 11572 11884 11612
rect 11924 11572 11925 11612
rect 11883 11563 11925 11572
rect 8995 11528 9053 11529
rect 8995 11488 9004 11528
rect 9044 11488 9053 11528
rect 8995 11487 9053 11488
rect 10443 11528 10485 11537
rect 10443 11488 10444 11528
rect 10484 11488 10485 11528
rect 10443 11479 10485 11488
rect 14275 11528 14333 11529
rect 14275 11488 14284 11528
rect 14324 11488 14333 11528
rect 14275 11487 14333 11488
rect 576 11360 14400 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 14400 11360
rect 576 11296 14400 11320
rect 651 11192 693 11201
rect 651 11152 652 11192
rect 692 11152 693 11192
rect 651 11143 693 11152
rect 7171 11192 7229 11193
rect 7171 11152 7180 11192
rect 7220 11152 7229 11192
rect 7171 11151 7229 11152
rect 9859 11192 9917 11193
rect 9859 11152 9868 11192
rect 9908 11152 9917 11192
rect 9859 11151 9917 11152
rect 14283 11192 14325 11201
rect 14283 11152 14284 11192
rect 14324 11152 14325 11192
rect 14283 11143 14325 11152
rect 2187 11108 2229 11117
rect 2187 11068 2188 11108
rect 2228 11068 2229 11108
rect 2187 11059 2229 11068
rect 4779 11108 4821 11117
rect 4779 11068 4780 11108
rect 4820 11068 4821 11108
rect 4779 11059 4821 11068
rect 7467 11108 7509 11117
rect 7467 11068 7468 11108
rect 7508 11068 7509 11108
rect 7467 11059 7509 11068
rect 12259 11108 12317 11109
rect 12259 11068 12268 11108
rect 12308 11068 12317 11108
rect 12259 11067 12317 11068
rect 2563 11024 2621 11025
rect 2563 10984 2572 11024
rect 2612 10984 2621 11024
rect 2563 10983 2621 10984
rect 3427 11024 3485 11025
rect 3427 10984 3436 11024
rect 3476 10984 3485 11024
rect 3427 10983 3485 10984
rect 5155 11024 5213 11025
rect 5155 10984 5164 11024
rect 5204 10984 5213 11024
rect 5155 10983 5213 10984
rect 6019 11024 6077 11025
rect 6019 10984 6028 11024
rect 6068 10984 6077 11024
rect 6019 10983 6077 10984
rect 7843 11024 7901 11025
rect 7843 10984 7852 11024
rect 7892 10984 7901 11024
rect 7843 10983 7901 10984
rect 8707 11024 8765 11025
rect 8707 10984 8716 11024
rect 8756 10984 8765 11024
rect 8707 10983 8765 10984
rect 10051 11024 10109 11025
rect 10051 10984 10060 11024
rect 10100 10984 10109 11024
rect 10051 10983 10109 10984
rect 11587 11024 11645 11025
rect 11587 10984 11596 11024
rect 11636 10984 11645 11024
rect 11587 10983 11645 10984
rect 11779 11024 11837 11025
rect 11779 10984 11788 11024
rect 11828 10984 11837 11024
rect 11779 10983 11837 10984
rect 12067 11024 12125 11025
rect 12067 10984 12076 11024
rect 12116 10984 12125 11024
rect 12067 10983 12125 10984
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 4587 10940 4629 10949
rect 4587 10900 4588 10940
rect 4628 10900 4629 10940
rect 4587 10891 4629 10900
rect 14083 10940 14141 10941
rect 14083 10900 14092 10940
rect 14132 10900 14141 10940
rect 14083 10899 14141 10900
rect 10723 10772 10781 10773
rect 10723 10732 10732 10772
rect 10772 10732 10781 10772
rect 10723 10731 10781 10732
rect 10915 10772 10973 10773
rect 10915 10732 10924 10772
rect 10964 10732 10973 10772
rect 10915 10731 10973 10732
rect 576 10604 14400 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 14400 10604
rect 576 10540 14400 10564
rect 5259 10436 5301 10445
rect 5259 10396 5260 10436
rect 5300 10396 5301 10436
rect 5259 10387 5301 10396
rect 6315 10352 6357 10361
rect 6315 10312 6316 10352
rect 6356 10312 6357 10352
rect 6315 10303 6357 10312
rect 6891 10352 6933 10361
rect 6891 10312 6892 10352
rect 6932 10312 6933 10352
rect 6891 10303 6933 10312
rect 7275 10352 7317 10361
rect 7275 10312 7276 10352
rect 7316 10312 7317 10352
rect 7275 10303 7317 10312
rect 9283 10352 9341 10353
rect 9283 10312 9292 10352
rect 9332 10312 9341 10352
rect 9283 10311 9341 10312
rect 12363 10352 12405 10361
rect 12363 10312 12364 10352
rect 12404 10312 12405 10352
rect 12363 10303 12405 10312
rect 4483 10268 4541 10269
rect 4483 10228 4492 10268
rect 4532 10228 4541 10268
rect 4483 10227 4541 10228
rect 4963 10184 5021 10185
rect 4963 10144 4972 10184
rect 5012 10144 5021 10184
rect 4963 10143 5021 10144
rect 5923 10184 5981 10185
rect 5923 10144 5932 10184
rect 5972 10144 5981 10184
rect 5923 10143 5981 10144
rect 9003 10184 9045 10193
rect 9003 10144 9004 10184
rect 9044 10144 9045 10184
rect 9003 10135 9045 10144
rect 9195 10184 9237 10193
rect 9195 10144 9196 10184
rect 9236 10144 9237 10184
rect 9195 10135 9237 10144
rect 9291 10184 9333 10193
rect 9291 10144 9292 10184
rect 9332 10144 9333 10184
rect 9291 10135 9333 10144
rect 9579 10184 9621 10193
rect 9579 10144 9580 10184
rect 9620 10144 9621 10184
rect 9579 10135 9621 10144
rect 9771 10184 9813 10193
rect 9771 10144 9772 10184
rect 9812 10144 9813 10184
rect 9771 10135 9813 10144
rect 9859 10184 9917 10185
rect 9859 10144 9868 10184
rect 9908 10144 9917 10184
rect 9859 10143 9917 10144
rect 10155 10184 10197 10193
rect 10155 10144 10156 10184
rect 10196 10144 10197 10184
rect 10155 10135 10197 10144
rect 10251 10184 10293 10193
rect 10251 10144 10252 10184
rect 10292 10144 10293 10184
rect 10251 10135 10293 10144
rect 10347 10184 10389 10193
rect 10347 10144 10348 10184
rect 10388 10144 10389 10184
rect 10347 10135 10389 10144
rect 10731 10184 10773 10193
rect 10731 10144 10732 10184
rect 10772 10144 10773 10184
rect 10731 10135 10773 10144
rect 11395 10184 11453 10185
rect 11395 10144 11404 10184
rect 11444 10144 11453 10184
rect 11395 10143 11453 10144
rect 11779 10184 11837 10185
rect 11779 10144 11788 10184
rect 11828 10144 11837 10184
rect 11779 10143 11837 10144
rect 11875 10184 11933 10185
rect 11875 10144 11884 10184
rect 11924 10144 11933 10184
rect 11875 10143 11933 10144
rect 13411 10184 13469 10185
rect 13411 10144 13420 10184
rect 13460 10144 13469 10184
rect 13411 10143 13469 10144
rect 9675 10100 9717 10109
rect 9675 10060 9676 10100
rect 9716 10060 9717 10100
rect 9675 10051 9717 10060
rect 10051 10016 10109 10017
rect 10051 9976 10060 10016
rect 10100 9976 10109 10016
rect 10051 9975 10109 9976
rect 11595 10016 11637 10025
rect 11595 9976 11596 10016
rect 11636 9976 11637 10016
rect 11595 9967 11637 9976
rect 12739 10016 12797 10017
rect 12739 9976 12748 10016
rect 12788 9976 12797 10016
rect 12739 9975 12797 9976
rect 576 9848 14400 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 14400 9848
rect 576 9784 14400 9808
rect 11211 9596 11253 9605
rect 11211 9556 11212 9596
rect 11252 9556 11253 9596
rect 11211 9547 11253 9556
rect 12171 9596 12213 9605
rect 12171 9556 12172 9596
rect 12212 9556 12213 9596
rect 12171 9547 12213 9556
rect 3139 9512 3197 9513
rect 3139 9472 3148 9512
rect 3188 9472 3197 9512
rect 3139 9471 3197 9472
rect 3235 9512 3293 9513
rect 3235 9472 3244 9512
rect 3284 9472 3293 9512
rect 3235 9471 3293 9472
rect 5259 9512 5301 9521
rect 5259 9472 5260 9512
rect 5300 9472 5301 9512
rect 5259 9463 5301 9472
rect 5451 9512 5493 9521
rect 5451 9472 5452 9512
rect 5492 9472 5493 9512
rect 5451 9463 5493 9472
rect 5643 9512 5685 9521
rect 5643 9472 5644 9512
rect 5684 9472 5685 9512
rect 5643 9463 5685 9472
rect 6019 9512 6077 9513
rect 6019 9472 6028 9512
rect 6068 9472 6077 9512
rect 6019 9471 6077 9472
rect 6883 9512 6941 9513
rect 6883 9472 6892 9512
rect 6932 9472 6941 9512
rect 6883 9471 6941 9472
rect 8131 9512 8189 9513
rect 8131 9472 8140 9512
rect 8180 9472 8189 9512
rect 8131 9471 8189 9472
rect 8523 9512 8565 9521
rect 8523 9472 8524 9512
rect 8564 9472 8565 9512
rect 8523 9463 8565 9472
rect 8899 9512 8957 9513
rect 8899 9472 8908 9512
rect 8948 9472 8957 9512
rect 8899 9471 8957 9472
rect 9763 9512 9821 9513
rect 9763 9472 9772 9512
rect 9812 9472 9821 9512
rect 9763 9471 9821 9472
rect 11307 9512 11349 9521
rect 11307 9472 11308 9512
rect 11348 9472 11349 9512
rect 11307 9463 11349 9472
rect 11403 9512 11445 9521
rect 11403 9472 11404 9512
rect 11444 9472 11445 9512
rect 11403 9463 11445 9472
rect 11499 9512 11541 9521
rect 11499 9472 11500 9512
rect 11540 9472 11541 9512
rect 11499 9463 11541 9472
rect 11779 9512 11837 9513
rect 11779 9472 11788 9512
rect 11828 9472 11837 9512
rect 11779 9471 11837 9472
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 12651 9512 12693 9521
rect 12651 9472 12652 9512
rect 12692 9472 12693 9512
rect 12651 9463 12693 9472
rect 13315 9512 13373 9513
rect 13315 9472 13324 9512
rect 13364 9472 13373 9512
rect 13315 9471 13373 9472
rect 13515 9512 13557 9521
rect 13515 9472 13516 9512
rect 13556 9472 13557 9512
rect 13515 9463 13557 9472
rect 13707 9512 13749 9521
rect 13707 9472 13708 9512
rect 13748 9472 13749 9512
rect 13707 9463 13749 9472
rect 13795 9512 13853 9513
rect 13795 9472 13804 9512
rect 13844 9472 13853 9512
rect 13795 9471 13853 9472
rect 2947 9428 3005 9429
rect 2947 9388 2956 9428
rect 2996 9388 3005 9428
rect 2947 9387 3005 9388
rect 3723 9344 3765 9353
rect 3723 9304 3724 9344
rect 3764 9304 3765 9344
rect 3723 9295 3765 9304
rect 5451 9344 5493 9353
rect 5451 9304 5452 9344
rect 5492 9304 5493 9344
rect 5451 9295 5493 9304
rect 13995 9344 14037 9353
rect 13995 9304 13996 9344
rect 14036 9304 14037 9344
rect 13995 9295 14037 9304
rect 10915 9260 10973 9261
rect 10915 9220 10924 9260
rect 10964 9220 10973 9260
rect 10915 9219 10973 9220
rect 12451 9260 12509 9261
rect 12451 9220 12460 9260
rect 12500 9220 12509 9260
rect 12451 9219 12509 9220
rect 13515 9260 13557 9269
rect 13515 9220 13516 9260
rect 13556 9220 13557 9260
rect 13515 9211 13557 9220
rect 576 9092 14400 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 14400 9092
rect 576 9028 14400 9052
rect 5547 8924 5589 8933
rect 5547 8884 5548 8924
rect 5588 8884 5589 8924
rect 5547 8875 5589 8884
rect 9003 8840 9045 8849
rect 9003 8800 9004 8840
rect 9044 8800 9045 8840
rect 9003 8791 9045 8800
rect 9387 8840 9429 8849
rect 9387 8800 9388 8840
rect 9428 8800 9429 8840
rect 9387 8791 9429 8800
rect 10443 8840 10485 8849
rect 10443 8800 10444 8840
rect 10484 8800 10485 8840
rect 10443 8791 10485 8800
rect 3331 8672 3389 8673
rect 3331 8632 3340 8672
rect 3380 8632 3389 8672
rect 3331 8631 3389 8632
rect 4195 8672 4253 8673
rect 4195 8632 4204 8672
rect 4244 8632 4253 8672
rect 4195 8631 4253 8632
rect 5635 8672 5693 8673
rect 5635 8632 5644 8672
rect 5684 8632 5693 8672
rect 5635 8631 5693 8632
rect 6211 8672 6269 8673
rect 6211 8632 6220 8672
rect 6260 8632 6269 8672
rect 6211 8631 6269 8632
rect 7075 8672 7133 8673
rect 7075 8632 7084 8672
rect 7124 8632 7133 8672
rect 7075 8631 7133 8632
rect 9475 8672 9533 8673
rect 9475 8632 9484 8672
rect 9524 8632 9533 8672
rect 9475 8631 9533 8632
rect 10251 8672 10293 8681
rect 10251 8632 10252 8672
rect 10292 8632 10293 8672
rect 10251 8623 10293 8632
rect 10347 8672 10389 8681
rect 10347 8632 10348 8672
rect 10388 8632 10389 8672
rect 10347 8623 10389 8632
rect 10539 8672 10581 8681
rect 10539 8632 10540 8672
rect 10580 8632 10581 8672
rect 10539 8623 10581 8632
rect 10915 8672 10973 8673
rect 10915 8632 10924 8672
rect 10964 8632 10973 8672
rect 10915 8631 10973 8632
rect 11595 8672 11637 8681
rect 11595 8632 11596 8672
rect 11636 8632 11637 8672
rect 11595 8623 11637 8632
rect 11787 8672 11829 8681
rect 11787 8632 11788 8672
rect 11828 8632 11829 8672
rect 11787 8623 11829 8632
rect 12163 8672 12221 8673
rect 12163 8632 12172 8672
rect 12212 8632 12221 8672
rect 12163 8631 12221 8632
rect 13027 8672 13085 8673
rect 13027 8632 13036 8672
rect 13076 8632 13085 8672
rect 13027 8631 13085 8632
rect 14187 8672 14229 8681
rect 14187 8632 14188 8672
rect 14228 8632 14229 8672
rect 14187 8623 14229 8632
rect 2955 8588 2997 8597
rect 2955 8548 2956 8588
rect 2996 8548 2997 8588
rect 2955 8539 2997 8548
rect 5835 8588 5877 8597
rect 5835 8548 5836 8588
rect 5876 8548 5877 8588
rect 5835 8539 5877 8548
rect 5347 8504 5405 8505
rect 5347 8464 5356 8504
rect 5396 8464 5405 8504
rect 5347 8463 5405 8464
rect 8227 8504 8285 8505
rect 8227 8464 8236 8504
rect 8276 8464 8285 8504
rect 8227 8463 8285 8464
rect 576 8336 14400 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 14400 8336
rect 576 8272 14400 8296
rect 4875 8199 4917 8208
rect 3043 8168 3101 8169
rect 3043 8128 3052 8168
rect 3092 8128 3101 8168
rect 3043 8127 3101 8128
rect 3331 8168 3389 8169
rect 3331 8128 3340 8168
rect 3380 8128 3389 8168
rect 3331 8127 3389 8128
rect 3523 8168 3581 8169
rect 3523 8128 3532 8168
rect 3572 8128 3581 8168
rect 4875 8159 4876 8199
rect 4916 8159 4917 8199
rect 4875 8150 4917 8159
rect 5923 8168 5981 8169
rect 3523 8127 3581 8128
rect 5923 8128 5932 8168
rect 5972 8128 5981 8168
rect 5923 8127 5981 8128
rect 11115 8168 11157 8177
rect 11115 8128 11116 8168
rect 11156 8128 11157 8168
rect 11115 8119 11157 8128
rect 11875 8168 11933 8169
rect 11875 8128 11884 8168
rect 11924 8128 11933 8168
rect 11875 8127 11933 8128
rect 9091 8084 9149 8085
rect 9091 8044 9100 8084
rect 9140 8044 9149 8084
rect 9091 8043 9149 8044
rect 14283 8084 14325 8093
rect 14283 8044 14284 8084
rect 14324 8044 14325 8084
rect 14283 8035 14325 8044
rect 2851 8000 2909 8001
rect 2851 7960 2860 8000
rect 2900 7960 2909 8000
rect 2851 7959 2909 7960
rect 3235 8000 3293 8001
rect 3235 7960 3244 8000
rect 3284 7960 3293 8000
rect 3235 7959 3293 7960
rect 4195 8000 4253 8001
rect 4195 7960 4204 8000
rect 4244 7960 4253 8000
rect 4195 7959 4253 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4771 8000 4829 8001
rect 4771 7960 4780 8000
rect 4820 7960 4829 8000
rect 4771 7959 4829 7960
rect 5059 8000 5117 8001
rect 5059 7960 5068 8000
rect 5108 7960 5117 8000
rect 5059 7959 5117 7960
rect 6595 8000 6653 8001
rect 6595 7960 6604 8000
rect 6644 7960 6653 8000
rect 6595 7959 6653 7960
rect 7459 8000 7517 8001
rect 7459 7960 7468 8000
rect 7508 7960 7517 8000
rect 7459 7959 7517 7960
rect 7747 8000 7805 8001
rect 7747 7960 7756 8000
rect 7796 7960 7805 8000
rect 7747 7959 7805 7960
rect 8707 8000 8765 8001
rect 8707 7960 8716 8000
rect 8756 7960 8765 8000
rect 8707 7959 8765 7960
rect 9187 8000 9245 8001
rect 9187 7960 9196 8000
rect 9236 7960 9245 8000
rect 9187 7959 9245 7960
rect 9571 8000 9629 8001
rect 9571 7960 9580 8000
rect 9620 7960 9629 8000
rect 9571 7959 9629 7960
rect 10155 8000 10197 8009
rect 10155 7960 10156 8000
rect 10196 7960 10197 8000
rect 10155 7951 10197 7960
rect 10347 8000 10389 8009
rect 10347 7960 10348 8000
rect 10388 7960 10389 8000
rect 10347 7951 10389 7960
rect 11299 8000 11357 8001
rect 11299 7960 11308 8000
rect 11348 7960 11357 8000
rect 11299 7959 11357 7960
rect 11587 8000 11645 8001
rect 11587 7960 11596 8000
rect 11636 7960 11645 8000
rect 11587 7959 11645 7960
rect 13027 8000 13085 8001
rect 13027 7960 13036 8000
rect 13076 7960 13085 8000
rect 13027 7959 13085 7960
rect 13891 8000 13949 8001
rect 13891 7960 13900 8000
rect 13940 7960 13949 8000
rect 13891 7959 13949 7960
rect 1611 7832 1653 7841
rect 1611 7792 1612 7832
rect 1652 7792 1653 7832
rect 1611 7783 1653 7792
rect 4395 7832 4437 7841
rect 4395 7792 4396 7832
rect 4436 7792 4437 7832
rect 4395 7783 4437 7792
rect 6787 7832 6845 7833
rect 6787 7792 6796 7832
rect 6836 7792 6845 7832
rect 6787 7791 6845 7792
rect 2179 7748 2237 7749
rect 2179 7708 2188 7748
rect 2228 7708 2237 7748
rect 2179 7707 2237 7708
rect 5731 7748 5789 7749
rect 5731 7708 5740 7748
rect 5780 7708 5789 7748
rect 5731 7707 5789 7708
rect 8043 7748 8085 7757
rect 8043 7708 8044 7748
rect 8084 7708 8085 7748
rect 8043 7699 8085 7708
rect 10347 7748 10389 7757
rect 10347 7708 10348 7748
rect 10388 7708 10389 7748
rect 10347 7699 10389 7708
rect 576 7580 14400 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 14400 7580
rect 576 7516 14400 7540
rect 4963 7412 5021 7413
rect 4963 7372 4972 7412
rect 5012 7372 5021 7412
rect 4963 7371 5021 7372
rect 5827 7412 5885 7413
rect 5827 7372 5836 7412
rect 5876 7372 5885 7412
rect 5827 7371 5885 7372
rect 11787 7328 11829 7337
rect 11787 7288 11788 7328
rect 11828 7288 11829 7328
rect 11787 7279 11829 7288
rect 1131 7160 1173 7169
rect 1131 7120 1132 7160
rect 1172 7120 1173 7160
rect 1131 7111 1173 7120
rect 1507 7160 1565 7161
rect 1507 7120 1516 7160
rect 1556 7120 1565 7160
rect 1507 7119 1565 7120
rect 2371 7160 2429 7161
rect 2371 7120 2380 7160
rect 2420 7120 2429 7160
rect 2371 7119 2429 7120
rect 4771 7160 4829 7161
rect 4771 7120 4780 7160
rect 4820 7120 4829 7160
rect 4771 7119 4829 7120
rect 5635 7160 5693 7161
rect 5635 7120 5644 7160
rect 5684 7120 5693 7160
rect 5635 7119 5693 7120
rect 6499 7160 6557 7161
rect 6499 7120 6508 7160
rect 6548 7120 6557 7160
rect 6499 7119 6557 7120
rect 7363 7160 7421 7161
rect 7363 7120 7372 7160
rect 7412 7120 7421 7160
rect 7363 7119 7421 7120
rect 8515 7160 8573 7161
rect 8515 7120 8524 7160
rect 8564 7120 8573 7160
rect 8515 7119 8573 7120
rect 8707 7160 8765 7161
rect 8707 7120 8716 7160
rect 8756 7120 8765 7160
rect 8707 7119 8765 7120
rect 8907 7160 8949 7169
rect 8907 7120 8908 7160
rect 8948 7120 8949 7160
rect 8907 7111 8949 7120
rect 9571 7160 9629 7161
rect 9571 7120 9580 7160
rect 9620 7120 9629 7160
rect 9571 7119 9629 7120
rect 10435 7160 10493 7161
rect 10435 7120 10444 7160
rect 10484 7120 10493 7160
rect 10435 7119 10493 7120
rect 8811 7076 8853 7085
rect 8811 7036 8812 7076
rect 8852 7036 8853 7076
rect 8811 7027 8853 7036
rect 9195 7076 9237 7085
rect 9195 7036 9196 7076
rect 9236 7036 9237 7076
rect 9195 7027 9237 7036
rect 3523 6992 3581 6993
rect 3523 6952 3532 6992
rect 3572 6952 3581 6992
rect 3523 6951 3581 6952
rect 4099 6992 4157 6993
rect 4099 6952 4108 6992
rect 4148 6952 4157 6992
rect 4099 6951 4157 6952
rect 4963 6992 5021 6993
rect 4963 6952 4972 6992
rect 5012 6952 5021 6992
rect 4963 6951 5021 6952
rect 6691 6992 6749 6993
rect 6691 6952 6700 6992
rect 6740 6952 6749 6992
rect 6691 6951 6749 6952
rect 7843 6992 7901 6993
rect 7843 6952 7852 6992
rect 7892 6952 7901 6992
rect 7843 6951 7901 6952
rect 11587 6992 11645 6993
rect 11587 6952 11596 6992
rect 11636 6952 11645 6992
rect 11587 6951 11645 6952
rect 576 6824 14400 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 14400 6824
rect 576 6760 14400 6784
rect 5931 6656 5973 6665
rect 5931 6616 5932 6656
rect 5972 6616 5973 6656
rect 5931 6607 5973 6616
rect 9187 6656 9245 6657
rect 9187 6616 9196 6656
rect 9236 6616 9245 6656
rect 9187 6615 9245 6616
rect 10723 6656 10781 6657
rect 10723 6616 10732 6656
rect 10772 6616 10781 6656
rect 10723 6615 10781 6616
rect 2667 6488 2709 6497
rect 2667 6448 2668 6488
rect 2708 6448 2709 6488
rect 2667 6439 2709 6448
rect 3043 6488 3101 6489
rect 3043 6448 3052 6488
rect 3092 6448 3101 6488
rect 3043 6447 3101 6448
rect 3907 6488 3965 6489
rect 3907 6448 3916 6488
rect 3956 6448 3965 6488
rect 3907 6447 3965 6448
rect 5547 6488 5589 6497
rect 5547 6448 5548 6488
rect 5588 6448 5589 6488
rect 5547 6439 5589 6448
rect 5635 6488 5693 6489
rect 5635 6448 5644 6488
rect 5684 6448 5693 6488
rect 5635 6447 5693 6448
rect 6211 6488 6269 6489
rect 6211 6448 6220 6488
rect 6260 6448 6269 6488
rect 6211 6447 6269 6448
rect 6411 6488 6453 6497
rect 6411 6448 6412 6488
rect 6452 6448 6453 6488
rect 6411 6439 6453 6448
rect 6787 6488 6845 6489
rect 6787 6448 6796 6488
rect 6836 6448 6845 6488
rect 6787 6447 6845 6448
rect 7651 6488 7709 6489
rect 7651 6448 7660 6488
rect 7700 6448 7709 6488
rect 7651 6447 7709 6448
rect 9859 6488 9917 6489
rect 9859 6448 9868 6488
rect 9908 6448 9917 6488
rect 9859 6447 9917 6448
rect 11395 6488 11453 6489
rect 11395 6448 11404 6488
rect 11444 6448 11453 6488
rect 11395 6447 11453 6448
rect 12547 6488 12605 6489
rect 12547 6448 12556 6488
rect 12596 6448 12605 6488
rect 12547 6447 12605 6448
rect 5067 6320 5109 6329
rect 5067 6280 5068 6320
rect 5108 6280 5109 6320
rect 5067 6271 5109 6280
rect 10059 6320 10101 6329
rect 10059 6280 10060 6320
rect 10100 6280 10101 6320
rect 10059 6271 10101 6280
rect 12747 6320 12789 6329
rect 12747 6280 12748 6320
rect 12788 6280 12789 6320
rect 12747 6271 12789 6280
rect 6123 6236 6165 6245
rect 6123 6196 6124 6236
rect 6164 6196 6165 6236
rect 6123 6187 6165 6196
rect 8803 6236 8861 6237
rect 8803 6196 8812 6236
rect 8852 6196 8861 6236
rect 8803 6195 8861 6196
rect 11875 6236 11933 6237
rect 11875 6196 11884 6236
rect 11924 6196 11933 6236
rect 11875 6195 11933 6196
rect 576 6068 14400 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 14400 6068
rect 576 6004 14400 6028
rect 4491 5900 4533 5909
rect 4491 5860 4492 5900
rect 4532 5860 4533 5900
rect 4491 5851 4533 5860
rect 5163 5900 5205 5909
rect 5163 5860 5164 5900
rect 5204 5860 5205 5900
rect 5163 5851 5205 5860
rect 6219 5900 6261 5909
rect 6219 5860 6220 5900
rect 6260 5860 6261 5900
rect 6219 5851 6261 5860
rect 8515 5900 8573 5901
rect 8515 5860 8524 5900
rect 8564 5860 8573 5900
rect 8515 5859 8573 5860
rect 9379 5900 9437 5901
rect 9379 5860 9388 5900
rect 9428 5860 9437 5900
rect 9379 5859 9437 5860
rect 1419 5816 1461 5825
rect 1419 5776 1420 5816
rect 1460 5776 1461 5816
rect 1419 5767 1461 5776
rect 3147 5816 3189 5825
rect 3147 5776 3148 5816
rect 3188 5776 3189 5816
rect 3147 5767 3189 5776
rect 4483 5648 4541 5649
rect 4483 5608 4492 5648
rect 4532 5608 4541 5648
rect 4483 5607 4541 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 4771 5648 4829 5649
rect 4771 5608 4780 5648
rect 4820 5608 4829 5648
rect 4771 5607 4829 5608
rect 4971 5648 5013 5657
rect 4971 5608 4972 5648
rect 5012 5608 5013 5648
rect 4971 5599 5013 5608
rect 5163 5648 5205 5657
rect 5163 5608 5164 5648
rect 5204 5608 5205 5648
rect 5163 5599 5205 5608
rect 5635 5648 5693 5649
rect 5635 5608 5644 5648
rect 5684 5608 5693 5648
rect 5635 5607 5693 5608
rect 5923 5648 5981 5649
rect 5923 5608 5932 5648
rect 5972 5608 5981 5648
rect 5923 5607 5981 5608
rect 6411 5648 6453 5657
rect 6411 5608 6412 5648
rect 6452 5608 6453 5648
rect 6411 5599 6453 5608
rect 6507 5648 6549 5657
rect 6507 5608 6508 5648
rect 6548 5608 6549 5648
rect 6507 5599 6549 5608
rect 6787 5648 6845 5649
rect 6787 5608 6796 5648
rect 6836 5608 6845 5648
rect 6787 5607 6845 5608
rect 7075 5648 7133 5649
rect 7075 5608 7084 5648
rect 7124 5608 7133 5648
rect 7075 5607 7133 5608
rect 7267 5648 7325 5649
rect 7267 5608 7276 5648
rect 7316 5608 7325 5648
rect 7267 5607 7325 5608
rect 7459 5648 7517 5649
rect 7459 5608 7468 5648
rect 7508 5608 7517 5648
rect 7459 5607 7517 5608
rect 8035 5648 8093 5649
rect 8035 5608 8044 5648
rect 8084 5608 8093 5648
rect 8035 5607 8093 5608
rect 8139 5648 8181 5657
rect 8139 5608 8140 5648
rect 8180 5608 8181 5648
rect 8139 5599 8181 5608
rect 8331 5648 8373 5657
rect 8331 5608 8332 5648
rect 8372 5608 8373 5648
rect 8331 5599 8373 5608
rect 9187 5648 9245 5649
rect 9187 5608 9196 5648
rect 9236 5608 9245 5648
rect 9187 5607 9245 5608
rect 10051 5648 10109 5649
rect 10051 5608 10060 5648
rect 10100 5608 10109 5648
rect 10051 5607 10109 5608
rect 10915 5648 10973 5649
rect 10915 5608 10924 5648
rect 10964 5608 10973 5648
rect 10915 5607 10973 5608
rect 11779 5648 11837 5649
rect 11779 5608 11788 5648
rect 11828 5608 11837 5648
rect 11779 5607 11837 5608
rect 5443 5564 5501 5565
rect 5443 5524 5452 5564
rect 5492 5524 5501 5564
rect 5443 5523 5501 5524
rect 6307 5564 6365 5565
rect 6307 5524 6316 5564
rect 6356 5524 6365 5564
rect 6307 5523 6365 5524
rect 10539 5564 10581 5573
rect 10539 5524 10540 5564
rect 10580 5524 10581 5564
rect 10539 5515 10581 5524
rect 6211 5480 6269 5481
rect 6211 5440 6220 5480
rect 6260 5440 6269 5480
rect 6211 5439 6269 5440
rect 7083 5480 7125 5489
rect 7083 5440 7084 5480
rect 7124 5440 7125 5480
rect 7083 5431 7125 5440
rect 8227 5480 8285 5481
rect 8227 5440 8236 5480
rect 8276 5440 8285 5480
rect 8227 5439 8285 5440
rect 12931 5480 12989 5481
rect 12931 5440 12940 5480
rect 12980 5440 12989 5480
rect 12931 5439 12989 5440
rect 576 5312 14400 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 14400 5312
rect 576 5248 14400 5272
rect 5355 5148 5397 5157
rect 5355 5108 5356 5148
rect 5396 5108 5397 5148
rect 5355 5099 5397 5108
rect 6019 5144 6077 5145
rect 6019 5104 6028 5144
rect 6068 5104 6077 5144
rect 6019 5103 6077 5104
rect 6603 5144 6645 5153
rect 6603 5104 6604 5144
rect 6644 5104 6645 5144
rect 6603 5095 6645 5104
rect 3811 5060 3869 5061
rect 3811 5020 3820 5060
rect 3860 5020 3869 5060
rect 3811 5019 3869 5020
rect 6987 5060 7029 5069
rect 6987 5020 6988 5060
rect 7028 5020 7029 5060
rect 6987 5011 7029 5020
rect 7851 5060 7893 5069
rect 7851 5020 7852 5060
rect 7892 5020 7893 5060
rect 7851 5011 7893 5020
rect 11883 5060 11925 5069
rect 11883 5020 11884 5060
rect 11924 5020 11925 5060
rect 11883 5011 11925 5020
rect 939 4976 981 4985
rect 939 4936 940 4976
rect 980 4936 981 4976
rect 939 4927 981 4936
rect 1315 4976 1373 4977
rect 1315 4936 1324 4976
rect 1364 4936 1373 4976
rect 1315 4935 1373 4936
rect 2179 4976 2237 4977
rect 2179 4936 2188 4976
rect 2228 4936 2237 4976
rect 2179 4935 2237 4936
rect 3427 4976 3485 4977
rect 3427 4936 3436 4976
rect 3476 4936 3485 4976
rect 3427 4935 3485 4936
rect 3907 4976 3965 4977
rect 3907 4936 3916 4976
rect 3956 4936 3965 4976
rect 3907 4935 3965 4936
rect 4291 4976 4349 4977
rect 4291 4936 4300 4976
rect 4340 4936 4349 4976
rect 4291 4935 4349 4936
rect 5155 4976 5213 4977
rect 5155 4936 5164 4976
rect 5204 4936 5213 4976
rect 5155 4935 5213 4936
rect 5443 4976 5501 4977
rect 5443 4936 5452 4976
rect 5492 4936 5501 4976
rect 5443 4935 5501 4936
rect 5547 4976 5589 4985
rect 5547 4936 5548 4976
rect 5588 4936 5589 4976
rect 5547 4927 5589 4936
rect 6115 4976 6173 4977
rect 6115 4936 6124 4976
rect 6164 4936 6173 4976
rect 6115 4935 6173 4936
rect 6507 4976 6549 4985
rect 6507 4936 6508 4976
rect 6548 4936 6549 4976
rect 6507 4927 6549 4936
rect 6699 4976 6741 4985
rect 6699 4936 6700 4976
rect 6740 4936 6741 4976
rect 6699 4927 6741 4936
rect 6795 4976 6837 4985
rect 6795 4936 6796 4976
rect 6836 4936 6837 4976
rect 6795 4927 6837 4936
rect 7651 4976 7709 4977
rect 7651 4936 7660 4976
rect 7700 4936 7709 4976
rect 7651 4935 7709 4936
rect 8227 4976 8285 4977
rect 8227 4936 8236 4976
rect 8276 4936 8285 4976
rect 8227 4935 8285 4936
rect 9091 4976 9149 4977
rect 9091 4936 9100 4976
rect 9140 4936 9149 4976
rect 9091 4935 9149 4936
rect 10635 4976 10677 4985
rect 10635 4936 10636 4976
rect 10676 4936 10677 4976
rect 10635 4927 10677 4936
rect 11491 4976 11549 4977
rect 11491 4936 11500 4976
rect 11540 4936 11549 4976
rect 11491 4935 11549 4936
rect 12259 4976 12317 4977
rect 12259 4936 12268 4976
rect 12308 4936 12317 4976
rect 12259 4935 12317 4936
rect 13123 4976 13181 4977
rect 13123 4936 13132 4976
rect 13172 4936 13181 4976
rect 13123 4935 13181 4936
rect 10251 4892 10293 4901
rect 10251 4852 10252 4892
rect 10292 4852 10293 4892
rect 10251 4843 10293 4852
rect 5835 4808 5877 4817
rect 5835 4768 5836 4808
rect 5876 4768 5877 4808
rect 5835 4759 5877 4768
rect 10827 4808 10869 4817
rect 10827 4768 10828 4808
rect 10868 4768 10869 4808
rect 10827 4759 10869 4768
rect 4483 4724 4541 4725
rect 4483 4684 4492 4724
rect 4532 4684 4541 4724
rect 4483 4683 4541 4684
rect 6307 4724 6365 4725
rect 6307 4684 6316 4724
rect 6356 4684 6365 4724
rect 6307 4683 6365 4684
rect 11019 4724 11061 4733
rect 11019 4684 11020 4724
rect 11060 4684 11061 4724
rect 11019 4675 11061 4684
rect 14275 4724 14333 4725
rect 14275 4684 14284 4724
rect 14324 4684 14333 4724
rect 14275 4683 14333 4684
rect 576 4556 14400 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 14400 4556
rect 576 4492 14400 4516
rect 1611 4388 1653 4397
rect 1611 4348 1612 4388
rect 1652 4348 1653 4388
rect 1611 4339 1653 4348
rect 7563 4388 7605 4397
rect 7563 4348 7564 4388
rect 7604 4348 7605 4388
rect 7563 4339 7605 4348
rect 10531 4388 10589 4389
rect 10531 4348 10540 4388
rect 10580 4348 10589 4388
rect 10531 4347 10589 4348
rect 11395 4388 11453 4389
rect 11395 4348 11404 4388
rect 11444 4348 11453 4388
rect 11395 4347 11453 4348
rect 2091 4304 2133 4313
rect 2091 4264 2092 4304
rect 2132 4264 2133 4304
rect 2091 4255 2133 4264
rect 2475 4304 2517 4313
rect 2475 4264 2476 4304
rect 2516 4264 2517 4304
rect 2475 4255 2517 4264
rect 3627 4304 3669 4313
rect 3627 4264 3628 4304
rect 3668 4264 3669 4304
rect 3627 4255 3669 4264
rect 8331 4304 8373 4313
rect 8331 4264 8332 4304
rect 8372 4264 8373 4304
rect 8331 4255 8373 4264
rect 14083 4220 14141 4221
rect 14083 4180 14092 4220
rect 14132 4180 14141 4220
rect 14083 4179 14141 4180
rect 1699 4136 1757 4137
rect 1699 4096 1708 4136
rect 1748 4096 1757 4136
rect 1699 4095 1757 4096
rect 2667 4136 2709 4145
rect 2667 4096 2668 4136
rect 2708 4096 2709 4136
rect 2667 4087 2709 4096
rect 3331 4136 3389 4137
rect 3331 4096 3340 4136
rect 3380 4096 3389 4136
rect 3331 4095 3389 4096
rect 4003 4136 4061 4137
rect 4003 4096 4012 4136
rect 4052 4096 4061 4136
rect 4003 4095 4061 4096
rect 4875 4136 4917 4145
rect 4875 4096 4876 4136
rect 4916 4096 4917 4136
rect 4875 4087 4917 4096
rect 6115 4136 6173 4137
rect 6115 4096 6124 4136
rect 6164 4096 6173 4136
rect 6115 4095 6173 4096
rect 6499 4136 6557 4137
rect 6499 4096 6508 4136
rect 6548 4096 6557 4136
rect 6499 4095 6557 4096
rect 7275 4136 7317 4145
rect 7275 4096 7276 4136
rect 7316 4096 7317 4136
rect 7275 4087 7317 4096
rect 7363 4136 7421 4137
rect 7363 4096 7372 4136
rect 7412 4096 7421 4136
rect 7363 4095 7421 4096
rect 7939 4136 7997 4137
rect 7939 4096 7948 4136
rect 7988 4096 7997 4136
rect 7939 4095 7997 4096
rect 8715 4136 8757 4145
rect 8715 4096 8716 4136
rect 8756 4096 8757 4136
rect 8715 4087 8757 4096
rect 8907 4136 8949 4145
rect 8907 4096 8908 4136
rect 8948 4096 8949 4136
rect 8907 4087 8949 4096
rect 10051 4136 10109 4137
rect 10051 4096 10060 4136
rect 10100 4096 10109 4136
rect 10051 4095 10109 4096
rect 11203 4136 11261 4137
rect 11203 4096 11212 4136
rect 11252 4096 11261 4136
rect 11203 4095 11261 4096
rect 12067 4136 12125 4137
rect 12067 4096 12076 4136
rect 12116 4096 12125 4136
rect 12067 4095 12125 4096
rect 12931 4136 12989 4137
rect 12931 4096 12940 4136
rect 12980 4096 12989 4136
rect 12931 4095 12989 4096
rect 13795 4136 13853 4137
rect 13795 4096 13804 4136
rect 13844 4096 13853 4136
rect 13795 4095 13853 4096
rect 5451 4052 5493 4061
rect 5451 4012 5452 4052
rect 5492 4012 5493 4052
rect 5451 4003 5493 4012
rect 6403 3968 6461 3969
rect 6403 3928 6412 3968
rect 6452 3928 6461 3968
rect 6403 3927 6461 3928
rect 6691 3968 6749 3969
rect 6691 3928 6700 3968
rect 6740 3928 6749 3968
rect 6691 3927 6749 3928
rect 7843 3968 7901 3969
rect 7843 3928 7852 3968
rect 7892 3928 7901 3968
rect 7843 3927 7901 3928
rect 8131 3968 8189 3969
rect 8131 3928 8140 3968
rect 8180 3928 8189 3968
rect 8131 3927 8189 3928
rect 8811 3968 8853 3977
rect 8811 3928 8812 3968
rect 8852 3928 8853 3968
rect 8811 3919 8853 3928
rect 9379 3968 9437 3969
rect 9379 3928 9388 3968
rect 9428 3928 9437 3968
rect 9379 3927 9437 3928
rect 12259 3968 12317 3969
rect 12259 3928 12268 3968
rect 12308 3928 12317 3968
rect 12259 3927 12317 3928
rect 13123 3968 13181 3969
rect 13123 3928 13132 3968
rect 13172 3928 13181 3968
rect 13123 3927 13181 3928
rect 14283 3968 14325 3977
rect 14283 3928 14284 3968
rect 14324 3928 14325 3968
rect 14283 3919 14325 3928
rect 576 3800 14400 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 14400 3800
rect 576 3736 14400 3760
rect 6987 3690 7029 3699
rect 6987 3650 6988 3690
rect 7028 3650 7029 3690
rect 6987 3641 7029 3650
rect 5059 3632 5117 3633
rect 5059 3592 5068 3632
rect 5108 3592 5117 3632
rect 5059 3591 5117 3592
rect 10819 3632 10877 3633
rect 10819 3592 10828 3632
rect 10868 3592 10877 3632
rect 10819 3591 10877 3592
rect 11211 3632 11253 3641
rect 11211 3592 11212 3632
rect 11252 3592 11253 3632
rect 11211 3583 11253 3592
rect 2667 3548 2709 3557
rect 2667 3508 2668 3548
rect 2708 3508 2709 3548
rect 2667 3499 2709 3508
rect 6595 3548 6653 3549
rect 6595 3508 6604 3548
rect 6644 3508 6653 3548
rect 6595 3507 6653 3508
rect 8131 3548 8189 3549
rect 8131 3508 8140 3548
rect 8180 3508 8189 3548
rect 8131 3507 8189 3508
rect 11979 3548 12021 3557
rect 11979 3508 11980 3548
rect 12020 3508 12021 3548
rect 11979 3499 12021 3508
rect 3043 3464 3101 3465
rect 3043 3424 3052 3464
rect 3092 3424 3101 3464
rect 3043 3423 3101 3424
rect 3907 3464 3965 3465
rect 3907 3424 3916 3464
rect 3956 3424 3965 3464
rect 3907 3423 3965 3424
rect 5355 3464 5397 3473
rect 5355 3424 5356 3464
rect 5396 3424 5397 3464
rect 5355 3415 5397 3424
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5443 3422 5501 3423
rect 5443 3382 5452 3422
rect 5492 3382 5501 3422
rect 5547 3415 5589 3424
rect 5643 3464 5685 3473
rect 5643 3424 5644 3464
rect 5684 3424 5685 3464
rect 5643 3415 5685 3424
rect 6115 3464 6173 3465
rect 6115 3424 6124 3464
rect 6164 3424 6173 3464
rect 6115 3423 6173 3424
rect 6403 3464 6461 3465
rect 6403 3424 6412 3464
rect 6452 3424 6461 3464
rect 6403 3423 6461 3424
rect 7075 3464 7133 3465
rect 7075 3424 7084 3464
rect 7124 3424 7133 3464
rect 7075 3423 7133 3424
rect 7179 3464 7221 3473
rect 7179 3424 7180 3464
rect 7220 3424 7221 3464
rect 7179 3415 7221 3424
rect 7651 3464 7709 3465
rect 7651 3424 7660 3464
rect 7700 3424 7709 3464
rect 7651 3423 7709 3424
rect 7939 3464 7997 3465
rect 7939 3424 7948 3464
rect 7988 3424 7997 3464
rect 7939 3423 7997 3424
rect 8419 3464 8477 3465
rect 8419 3424 8428 3464
rect 8468 3424 8477 3464
rect 8419 3423 8477 3424
rect 10051 3464 10109 3465
rect 10051 3424 10060 3464
rect 10100 3424 10109 3464
rect 10051 3423 10109 3424
rect 10627 3464 10685 3465
rect 10627 3424 10636 3464
rect 10676 3424 10685 3464
rect 10627 3423 10685 3424
rect 10731 3464 10773 3473
rect 10731 3424 10732 3464
rect 10772 3424 10773 3464
rect 10731 3415 10773 3424
rect 10923 3464 10965 3473
rect 10923 3424 10924 3464
rect 10964 3424 10965 3464
rect 10923 3415 10965 3424
rect 11299 3464 11357 3465
rect 11299 3424 11308 3464
rect 11348 3424 11357 3464
rect 11299 3423 11357 3424
rect 11683 3464 11741 3465
rect 11683 3424 11692 3464
rect 11732 3424 11741 3464
rect 11683 3423 11741 3424
rect 11875 3464 11933 3465
rect 11875 3424 11884 3464
rect 11924 3424 11933 3464
rect 11875 3423 11933 3424
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 5443 3381 5501 3382
rect 9387 3380 9429 3389
rect 9387 3340 9388 3380
rect 9428 3340 9429 3380
rect 9387 3331 9429 3340
rect 5827 3296 5885 3297
rect 5827 3256 5836 3296
rect 5876 3256 5885 3296
rect 5827 3255 5885 3256
rect 7467 3296 7509 3305
rect 7467 3256 7468 3296
rect 7508 3256 7509 3296
rect 7467 3247 7509 3256
rect 10251 3296 10293 3305
rect 10251 3256 10252 3296
rect 10292 3256 10293 3296
rect 10251 3247 10293 3256
rect 9091 3212 9149 3213
rect 9091 3172 9100 3212
rect 9140 3172 9149 3212
rect 9091 3171 9149 3172
rect 576 3044 14400 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 14400 3044
rect 576 2980 14400 3004
rect 4387 2876 4445 2877
rect 4387 2836 4396 2876
rect 4436 2836 4445 2876
rect 4387 2835 4445 2836
rect 4779 2876 4821 2885
rect 4779 2836 4780 2876
rect 4820 2836 4821 2876
rect 4779 2827 4821 2836
rect 5251 2876 5309 2877
rect 5251 2836 5260 2876
rect 5300 2836 5309 2876
rect 5251 2835 5309 2836
rect 10819 2876 10877 2877
rect 10819 2836 10828 2876
rect 10868 2836 10877 2876
rect 10819 2835 10877 2836
rect 11011 2708 11069 2709
rect 11011 2668 11020 2708
rect 11060 2668 11069 2708
rect 11011 2667 11069 2668
rect 1995 2624 2037 2633
rect 1995 2584 1996 2624
rect 2036 2584 2037 2624
rect 1995 2575 2037 2584
rect 2371 2624 2429 2625
rect 2371 2584 2380 2624
rect 2420 2584 2429 2624
rect 2371 2583 2429 2584
rect 3235 2624 3293 2625
rect 3235 2584 3244 2624
rect 3284 2584 3293 2624
rect 3235 2583 3293 2584
rect 4771 2624 4829 2625
rect 4771 2584 4780 2624
rect 4820 2584 4829 2624
rect 4771 2583 4829 2584
rect 4971 2624 5013 2633
rect 4971 2584 4972 2624
rect 5012 2584 5013 2624
rect 4971 2575 5013 2584
rect 5059 2624 5117 2625
rect 5059 2584 5068 2624
rect 5108 2584 5117 2624
rect 5059 2583 5117 2584
rect 5923 2624 5981 2625
rect 5923 2584 5932 2624
rect 5972 2584 5981 2624
rect 5923 2583 5981 2584
rect 6115 2624 6173 2625
rect 6115 2584 6124 2624
rect 6164 2584 6173 2624
rect 6115 2583 6173 2584
rect 6987 2624 7029 2633
rect 6987 2584 6988 2624
rect 7028 2584 7029 2624
rect 6987 2575 7029 2584
rect 7083 2624 7125 2633
rect 7083 2584 7084 2624
rect 7124 2584 7125 2624
rect 7083 2575 7125 2584
rect 7555 2624 7613 2625
rect 7555 2584 7564 2624
rect 7604 2584 7613 2624
rect 7555 2583 7613 2584
rect 8427 2624 8469 2633
rect 8427 2584 8428 2624
rect 8468 2584 8469 2624
rect 8427 2575 8469 2584
rect 8803 2624 8861 2625
rect 8803 2584 8812 2624
rect 8852 2584 8861 2624
rect 8803 2583 8861 2584
rect 9667 2624 9725 2625
rect 9667 2584 9676 2624
rect 9716 2584 9725 2624
rect 9667 2583 9725 2584
rect 6795 2540 6837 2549
rect 6795 2500 6796 2540
rect 6836 2500 6837 2540
rect 6795 2491 6837 2500
rect 7171 2540 7229 2541
rect 7171 2500 7180 2540
rect 7220 2500 7229 2540
rect 7171 2499 7229 2500
rect 5251 2456 5309 2457
rect 5251 2416 5260 2456
rect 5300 2416 5309 2456
rect 5251 2415 5309 2416
rect 7267 2456 7325 2457
rect 7267 2416 7276 2456
rect 7316 2416 7325 2456
rect 7267 2415 7325 2416
rect 7371 2456 7413 2465
rect 7371 2416 7372 2456
rect 7412 2416 7413 2456
rect 7371 2407 7413 2416
rect 8227 2456 8285 2457
rect 8227 2416 8236 2456
rect 8276 2416 8285 2456
rect 8227 2415 8285 2416
rect 576 2288 14400 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 14400 2288
rect 576 2224 14400 2248
rect 5539 2120 5597 2121
rect 5539 2080 5548 2120
rect 5588 2080 5597 2120
rect 5539 2079 5597 2080
rect 5923 2120 5981 2121
rect 5923 2080 5932 2120
rect 5972 2080 5981 2120
rect 5923 2079 5981 2080
rect 10915 2120 10973 2121
rect 10915 2080 10924 2120
rect 10964 2080 10973 2120
rect 10915 2079 10973 2080
rect 8331 2036 8373 2045
rect 8331 1996 8332 2036
rect 8372 1996 8373 2036
rect 8331 1987 8373 1996
rect 8523 2036 8565 2045
rect 8523 1996 8524 2036
rect 8564 1996 8565 2036
rect 8523 1987 8565 1996
rect 3147 1952 3189 1961
rect 3147 1912 3148 1952
rect 3188 1912 3189 1952
rect 3147 1903 3189 1912
rect 3523 1952 3581 1953
rect 3523 1912 3532 1952
rect 3572 1912 3581 1952
rect 3523 1911 3581 1912
rect 4387 1952 4445 1953
rect 4387 1912 4396 1952
rect 4436 1912 4445 1952
rect 4387 1911 4445 1912
rect 7075 1952 7133 1953
rect 7075 1912 7084 1952
rect 7124 1912 7133 1952
rect 7075 1911 7133 1912
rect 7939 1952 7997 1953
rect 7939 1912 7948 1952
rect 7988 1912 7997 1952
rect 7939 1911 7997 1912
rect 8899 1952 8957 1953
rect 8899 1912 8908 1952
rect 8948 1912 8957 1952
rect 8899 1911 8957 1912
rect 9763 1952 9821 1953
rect 9763 1912 9772 1952
rect 9812 1912 9821 1952
rect 9763 1911 9821 1912
rect 576 1532 14400 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 14400 1532
rect 576 1468 14400 1492
rect 4099 1280 4157 1281
rect 4099 1240 4108 1280
rect 4148 1240 4157 1280
rect 4099 1239 4157 1240
rect 7083 1280 7125 1289
rect 7083 1240 7084 1280
rect 7124 1240 7125 1280
rect 7083 1231 7125 1240
rect 9387 1280 9429 1289
rect 9387 1240 9388 1280
rect 9428 1240 9429 1280
rect 9387 1231 9429 1240
rect 4963 1196 5021 1197
rect 4963 1156 4972 1196
rect 5012 1156 5021 1196
rect 4963 1155 5021 1156
rect 4771 1112 4829 1113
rect 4771 1072 4780 1112
rect 4820 1072 4829 1112
rect 4771 1071 4829 1072
rect 5251 1112 5309 1113
rect 5251 1072 5260 1112
rect 5300 1072 5309 1112
rect 5251 1071 5309 1072
rect 5355 1112 5397 1121
rect 5355 1072 5356 1112
rect 5396 1072 5397 1112
rect 5355 1063 5397 1072
rect 576 776 14400 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 14400 776
rect 576 712 14400 736
<< via1 >>
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 5260 13336 5300 13376
rect 6892 13336 6932 13376
rect 11212 13336 11252 13376
rect 7084 13168 7124 13208
rect 7180 13168 7220 13208
rect 7372 13168 7412 13208
rect 8236 13168 8276 13208
rect 8812 13168 8852 13208
rect 8908 13168 8948 13208
rect 9484 13168 9524 13208
rect 10156 13168 10196 13208
rect 10348 13168 10388 13208
rect 10540 13168 10580 13208
rect 10924 13168 10964 13208
rect 12364 13168 12404 13208
rect 9100 13084 9140 13124
rect 7276 13000 7316 13040
rect 7564 13000 7604 13040
rect 8812 13000 8852 13040
rect 10444 13000 10484 13040
rect 10732 13000 10772 13040
rect 11020 13000 11060 13040
rect 11692 13000 11732 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 7660 12664 7700 12704
rect 8428 12580 8468 12620
rect 3436 12496 3476 12536
rect 4780 12496 4820 12536
rect 4972 12496 5012 12536
rect 5260 12496 5300 12536
rect 5452 12496 5492 12536
rect 6124 12496 6164 12536
rect 7276 12496 7316 12536
rect 7468 12496 7508 12536
rect 7852 12496 7892 12536
rect 7948 12496 7988 12536
rect 9100 12496 9140 12536
rect 9964 12496 10004 12536
rect 10348 12496 10388 12536
rect 10732 12496 10772 12536
rect 11596 12496 11636 12536
rect 1132 12328 1172 12368
rect 2572 12328 2612 12368
rect 3724 12328 3764 12368
rect 6796 12328 6836 12368
rect 12940 12328 12980 12368
rect 2764 12244 2804 12284
rect 4108 12244 4148 12284
rect 5260 12244 5300 12284
rect 7276 12244 7316 12284
rect 9292 12244 9332 12284
rect 12748 12244 12788 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3052 11908 3092 11948
rect 5740 11908 5780 11948
rect 8716 11824 8756 11864
rect 1036 11656 1076 11696
rect 1900 11656 1940 11696
rect 3340 11656 3380 11696
rect 3724 11656 3764 11696
rect 4588 11656 4628 11696
rect 6316 11656 6356 11696
rect 6700 11656 6740 11696
rect 7564 11656 7604 11696
rect 9676 11656 9716 11696
rect 10060 11656 10100 11696
rect 10156 11656 10196 11696
rect 10828 11656 10868 11696
rect 11692 11656 11732 11696
rect 12268 11656 12308 11696
rect 13132 11656 13172 11696
rect 652 11572 692 11612
rect 11884 11572 11924 11612
rect 9004 11488 9044 11528
rect 10444 11488 10484 11528
rect 14284 11488 14324 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 652 11152 692 11192
rect 7180 11152 7220 11192
rect 9868 11152 9908 11192
rect 14284 11152 14324 11192
rect 2188 11068 2228 11108
rect 4780 11068 4820 11108
rect 7468 11068 7508 11108
rect 12268 11068 12308 11108
rect 2572 10984 2612 11024
rect 3436 10984 3476 11024
rect 5164 10984 5204 11024
rect 6028 10984 6068 11024
rect 7852 10984 7892 11024
rect 8716 10984 8756 11024
rect 10060 10984 10100 11024
rect 11596 10984 11636 11024
rect 11788 10984 11828 11024
rect 12076 10984 12116 11024
rect 844 10900 884 10940
rect 4588 10900 4628 10940
rect 14092 10900 14132 10940
rect 10732 10732 10772 10772
rect 10924 10732 10964 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 5260 10396 5300 10436
rect 6316 10312 6356 10352
rect 6892 10312 6932 10352
rect 7276 10312 7316 10352
rect 9292 10312 9332 10352
rect 12364 10312 12404 10352
rect 4492 10228 4532 10268
rect 4972 10144 5012 10184
rect 5932 10144 5972 10184
rect 9004 10144 9044 10184
rect 9196 10144 9236 10184
rect 9292 10144 9332 10184
rect 9580 10144 9620 10184
rect 9772 10144 9812 10184
rect 9868 10144 9908 10184
rect 10156 10144 10196 10184
rect 10252 10144 10292 10184
rect 10348 10144 10388 10184
rect 10732 10144 10772 10184
rect 11404 10144 11444 10184
rect 11788 10144 11828 10184
rect 11884 10144 11924 10184
rect 13420 10144 13460 10184
rect 9676 10060 9716 10100
rect 10060 9976 10100 10016
rect 11596 9976 11636 10016
rect 12748 9976 12788 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 11212 9556 11252 9596
rect 12172 9556 12212 9596
rect 3148 9472 3188 9512
rect 3244 9472 3284 9512
rect 5260 9472 5300 9512
rect 5452 9472 5492 9512
rect 5644 9472 5684 9512
rect 6028 9472 6068 9512
rect 6892 9472 6932 9512
rect 8140 9472 8180 9512
rect 8524 9472 8564 9512
rect 8908 9472 8948 9512
rect 9772 9472 9812 9512
rect 11308 9472 11348 9512
rect 11404 9472 11444 9512
rect 11500 9472 11540 9512
rect 11788 9472 11828 9512
rect 12076 9472 12116 9512
rect 12652 9472 12692 9512
rect 13324 9472 13364 9512
rect 13516 9472 13556 9512
rect 13708 9472 13748 9512
rect 13804 9472 13844 9512
rect 2956 9388 2996 9428
rect 3724 9304 3764 9344
rect 5452 9304 5492 9344
rect 13996 9304 14036 9344
rect 10924 9220 10964 9260
rect 12460 9220 12500 9260
rect 13516 9220 13556 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 5548 8884 5588 8924
rect 9004 8800 9044 8840
rect 9388 8800 9428 8840
rect 10444 8800 10484 8840
rect 3340 8632 3380 8672
rect 4204 8632 4244 8672
rect 5644 8632 5684 8672
rect 6220 8632 6260 8672
rect 7084 8632 7124 8672
rect 9484 8632 9524 8672
rect 10252 8632 10292 8672
rect 10348 8632 10388 8672
rect 10540 8632 10580 8672
rect 10924 8632 10964 8672
rect 11596 8632 11636 8672
rect 11788 8632 11828 8672
rect 12172 8632 12212 8672
rect 13036 8632 13076 8672
rect 14188 8632 14228 8672
rect 2956 8548 2996 8588
rect 5836 8548 5876 8588
rect 5356 8464 5396 8504
rect 8236 8464 8276 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3052 8128 3092 8168
rect 3340 8128 3380 8168
rect 3532 8128 3572 8168
rect 4876 8159 4916 8199
rect 5932 8128 5972 8168
rect 11116 8128 11156 8168
rect 11884 8128 11924 8168
rect 9100 8044 9140 8084
rect 14284 8044 14324 8084
rect 2860 7960 2900 8000
rect 3244 7960 3284 8000
rect 4204 7960 4244 8000
rect 4684 7960 4724 8000
rect 4780 7960 4820 8000
rect 5068 7960 5108 8000
rect 6604 7960 6644 8000
rect 7468 7960 7508 8000
rect 7756 7960 7796 8000
rect 8716 7960 8756 8000
rect 9196 7960 9236 8000
rect 9580 7960 9620 8000
rect 10156 7960 10196 8000
rect 10348 7960 10388 8000
rect 11308 7960 11348 8000
rect 11596 7960 11636 8000
rect 13036 7960 13076 8000
rect 13900 7960 13940 8000
rect 1612 7792 1652 7832
rect 4396 7792 4436 7832
rect 6796 7792 6836 7832
rect 2188 7708 2228 7748
rect 5740 7708 5780 7748
rect 8044 7708 8084 7748
rect 10348 7708 10388 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4972 7372 5012 7412
rect 5836 7372 5876 7412
rect 11788 7288 11828 7328
rect 1132 7120 1172 7160
rect 1516 7120 1556 7160
rect 2380 7120 2420 7160
rect 4780 7120 4820 7160
rect 5644 7120 5684 7160
rect 6508 7120 6548 7160
rect 7372 7120 7412 7160
rect 8524 7120 8564 7160
rect 8716 7120 8756 7160
rect 8908 7120 8948 7160
rect 9580 7120 9620 7160
rect 10444 7120 10484 7160
rect 8812 7036 8852 7076
rect 9196 7036 9236 7076
rect 3532 6952 3572 6992
rect 4108 6952 4148 6992
rect 4972 6952 5012 6992
rect 6700 6952 6740 6992
rect 7852 6952 7892 6992
rect 11596 6952 11636 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 5932 6616 5972 6656
rect 9196 6616 9236 6656
rect 10732 6616 10772 6656
rect 2668 6448 2708 6488
rect 3052 6448 3092 6488
rect 3916 6448 3956 6488
rect 5548 6448 5588 6488
rect 5644 6448 5684 6488
rect 6220 6448 6260 6488
rect 6412 6448 6452 6488
rect 6796 6448 6836 6488
rect 7660 6448 7700 6488
rect 9868 6448 9908 6488
rect 11404 6448 11444 6488
rect 12556 6448 12596 6488
rect 5068 6280 5108 6320
rect 10060 6280 10100 6320
rect 12748 6280 12788 6320
rect 6124 6196 6164 6236
rect 8812 6196 8852 6236
rect 11884 6196 11924 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4492 5860 4532 5900
rect 5164 5860 5204 5900
rect 6220 5860 6260 5900
rect 8524 5860 8564 5900
rect 9388 5860 9428 5900
rect 1420 5776 1460 5816
rect 3148 5776 3188 5816
rect 4492 5608 4532 5648
rect 4684 5608 4724 5648
rect 4780 5608 4820 5648
rect 4972 5608 5012 5648
rect 5164 5608 5204 5648
rect 5644 5608 5684 5648
rect 5932 5608 5972 5648
rect 6412 5608 6452 5648
rect 6508 5608 6548 5648
rect 6796 5608 6836 5648
rect 7084 5608 7124 5648
rect 7276 5608 7316 5648
rect 7468 5608 7508 5648
rect 8044 5608 8084 5648
rect 8140 5608 8180 5648
rect 8332 5608 8372 5648
rect 9196 5608 9236 5648
rect 10060 5608 10100 5648
rect 10924 5608 10964 5648
rect 11788 5608 11828 5648
rect 5452 5524 5492 5564
rect 6316 5524 6356 5564
rect 10540 5524 10580 5564
rect 6220 5440 6260 5480
rect 7084 5440 7124 5480
rect 8236 5440 8276 5480
rect 12940 5440 12980 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 5356 5108 5396 5148
rect 6028 5104 6068 5144
rect 6604 5104 6644 5144
rect 3820 5020 3860 5060
rect 6988 5020 7028 5060
rect 7852 5020 7892 5060
rect 11884 5020 11924 5060
rect 940 4936 980 4976
rect 1324 4936 1364 4976
rect 2188 4936 2228 4976
rect 3436 4936 3476 4976
rect 3916 4936 3956 4976
rect 4300 4936 4340 4976
rect 5164 4936 5204 4976
rect 5452 4936 5492 4976
rect 5548 4936 5588 4976
rect 6124 4936 6164 4976
rect 6508 4936 6548 4976
rect 6700 4936 6740 4976
rect 6796 4936 6836 4976
rect 7660 4936 7700 4976
rect 8236 4936 8276 4976
rect 9100 4936 9140 4976
rect 10636 4936 10676 4976
rect 11500 4936 11540 4976
rect 12268 4936 12308 4976
rect 13132 4936 13172 4976
rect 10252 4852 10292 4892
rect 5836 4768 5876 4808
rect 10828 4768 10868 4808
rect 4492 4684 4532 4724
rect 6316 4684 6356 4724
rect 11020 4684 11060 4724
rect 14284 4684 14324 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 1612 4348 1652 4388
rect 7564 4348 7604 4388
rect 10540 4348 10580 4388
rect 11404 4348 11444 4388
rect 2092 4264 2132 4304
rect 2476 4264 2516 4304
rect 3628 4264 3668 4304
rect 8332 4264 8372 4304
rect 14092 4180 14132 4220
rect 1708 4096 1748 4136
rect 2668 4096 2708 4136
rect 3340 4096 3380 4136
rect 4012 4096 4052 4136
rect 4876 4096 4916 4136
rect 6124 4096 6164 4136
rect 6508 4096 6548 4136
rect 7276 4096 7316 4136
rect 7372 4096 7412 4136
rect 7948 4096 7988 4136
rect 8716 4096 8756 4136
rect 8908 4096 8948 4136
rect 10060 4096 10100 4136
rect 11212 4096 11252 4136
rect 12076 4096 12116 4136
rect 12940 4096 12980 4136
rect 13804 4096 13844 4136
rect 5452 4012 5492 4052
rect 6412 3928 6452 3968
rect 6700 3928 6740 3968
rect 7852 3928 7892 3968
rect 8140 3928 8180 3968
rect 8812 3928 8852 3968
rect 9388 3928 9428 3968
rect 12268 3928 12308 3968
rect 13132 3928 13172 3968
rect 14284 3928 14324 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 6988 3650 7028 3690
rect 5068 3592 5108 3632
rect 10828 3592 10868 3632
rect 11212 3592 11252 3632
rect 2668 3508 2708 3548
rect 6604 3508 6644 3548
rect 8140 3508 8180 3548
rect 11980 3508 12020 3548
rect 3052 3424 3092 3464
rect 3916 3424 3956 3464
rect 5356 3424 5396 3464
rect 5548 3424 5588 3464
rect 5452 3382 5492 3422
rect 5644 3424 5684 3464
rect 6124 3424 6164 3464
rect 6412 3424 6452 3464
rect 7084 3424 7124 3464
rect 7180 3424 7220 3464
rect 7660 3424 7700 3464
rect 7948 3424 7988 3464
rect 8428 3424 8468 3464
rect 10060 3424 10100 3464
rect 10636 3424 10676 3464
rect 10732 3424 10772 3464
rect 10924 3424 10964 3464
rect 11308 3424 11348 3464
rect 11692 3424 11732 3464
rect 11884 3424 11924 3464
rect 12076 3424 12116 3464
rect 9388 3340 9428 3380
rect 5836 3256 5876 3296
rect 7468 3256 7508 3296
rect 10252 3256 10292 3296
rect 9100 3172 9140 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 4396 2836 4436 2876
rect 4780 2836 4820 2876
rect 5260 2836 5300 2876
rect 10828 2836 10868 2876
rect 11020 2668 11060 2708
rect 1996 2584 2036 2624
rect 2380 2584 2420 2624
rect 3244 2584 3284 2624
rect 4780 2584 4820 2624
rect 4972 2584 5012 2624
rect 5068 2584 5108 2624
rect 5932 2584 5972 2624
rect 6124 2584 6164 2624
rect 6988 2584 7028 2624
rect 7084 2584 7124 2624
rect 7564 2584 7604 2624
rect 8428 2584 8468 2624
rect 8812 2584 8852 2624
rect 9676 2584 9716 2624
rect 6796 2500 6836 2540
rect 7180 2500 7220 2540
rect 5260 2416 5300 2456
rect 7276 2416 7316 2456
rect 7372 2416 7412 2456
rect 8236 2416 8276 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 5548 2080 5588 2120
rect 5932 2080 5972 2120
rect 10924 2080 10964 2120
rect 8332 1996 8372 2036
rect 8524 1996 8564 2036
rect 3148 1912 3188 1952
rect 3532 1912 3572 1952
rect 4396 1912 4436 1952
rect 7084 1912 7124 1952
rect 7948 1912 7988 1952
rect 8908 1912 8948 1952
rect 9772 1912 9812 1952
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 4108 1240 4148 1280
rect 7084 1240 7124 1280
rect 9388 1240 9428 1280
rect 4972 1156 5012 1196
rect 4780 1072 4820 1112
rect 5260 1072 5300 1112
rect 5356 1072 5396 1112
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
<< metal2 >>
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 5260 13376 5300 13385
rect 5164 13336 5260 13376
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 3436 12536 3476 12545
rect 2956 12496 3436 12536
rect 1132 12368 1172 12377
rect 1036 12328 1132 12368
rect 1036 11696 1076 12328
rect 1132 12319 1172 12328
rect 2572 12368 2612 12377
rect 2187 12284 2229 12293
rect 2187 12244 2188 12284
rect 2228 12244 2229 12284
rect 2187 12235 2229 12244
rect 1036 11647 1076 11656
rect 1900 11696 1940 11705
rect 652 11612 692 11621
rect 652 11192 692 11572
rect 652 11143 692 11152
rect 843 11192 885 11201
rect 843 11152 844 11192
rect 884 11152 885 11192
rect 843 11143 885 11152
rect 844 10940 884 11143
rect 1900 11033 1940 11656
rect 2188 11108 2228 12235
rect 2188 11059 2228 11068
rect 1899 11024 1941 11033
rect 1899 10984 1900 11024
rect 1940 10984 1941 11024
rect 1899 10975 1941 10984
rect 2572 11024 2612 12328
rect 2763 12284 2805 12293
rect 2763 12244 2764 12284
rect 2804 12244 2805 12284
rect 2763 12235 2805 12244
rect 2764 12150 2804 12235
rect 2956 11948 2996 12496
rect 3436 12487 3476 12496
rect 4107 12536 4149 12545
rect 4107 12496 4108 12536
rect 4148 12496 4149 12536
rect 4107 12487 4149 12496
rect 4780 12536 4820 12545
rect 4971 12536 5013 12545
rect 4820 12496 4916 12536
rect 4780 12487 4820 12496
rect 3724 12368 3764 12377
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 3052 11948 3092 11957
rect 2956 11908 3052 11948
rect 3052 11899 3092 11908
rect 3339 11696 3381 11705
rect 3339 11656 3340 11696
rect 3380 11656 3381 11696
rect 3339 11647 3381 11656
rect 3724 11696 3764 12328
rect 4108 12284 4148 12487
rect 4108 11705 4148 12244
rect 4779 12284 4821 12293
rect 4779 12244 4780 12284
rect 4820 12244 4821 12284
rect 4779 12235 4821 12244
rect 3724 11647 3764 11656
rect 4107 11696 4149 11705
rect 4588 11696 4628 11705
rect 4107 11656 4108 11696
rect 4148 11656 4149 11696
rect 4107 11647 4149 11656
rect 4204 11656 4588 11696
rect 3340 11562 3380 11647
rect 4204 11033 4244 11656
rect 4588 11647 4628 11656
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4780 11108 4820 12235
rect 4780 11059 4820 11068
rect 2572 10975 2612 10984
rect 3435 11024 3477 11033
rect 3435 10984 3436 11024
rect 3476 10984 3477 11024
rect 3435 10975 3477 10984
rect 4203 11024 4245 11033
rect 4203 10984 4204 11024
rect 4244 10984 4245 11024
rect 4203 10975 4245 10984
rect 4491 11024 4533 11033
rect 4491 10984 4492 11024
rect 4532 10984 4533 11024
rect 4491 10975 4533 10984
rect 844 10891 884 10900
rect 3436 10890 3476 10975
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3148 9512 3188 9521
rect 2956 9428 2996 9437
rect 2860 9388 2956 9428
rect 2860 8000 2900 9388
rect 2956 9379 2996 9388
rect 3148 9260 3188 9472
rect 3244 9512 3284 9521
rect 3284 9472 3572 9512
rect 3244 9463 3284 9472
rect 2956 9220 3188 9260
rect 2956 8924 2996 9220
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 2956 8884 3188 8924
rect 2956 8588 2996 8597
rect 2956 8168 2996 8548
rect 3052 8168 3092 8177
rect 2956 8128 3052 8168
rect 3148 8168 3188 8884
rect 3339 8672 3381 8681
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 3340 8538 3380 8623
rect 3340 8168 3380 8177
rect 3148 8128 3340 8168
rect 3052 8119 3092 8128
rect 2860 7951 2900 7960
rect 3243 8000 3285 8009
rect 3243 7960 3244 8000
rect 3284 7960 3285 8000
rect 3243 7951 3285 7960
rect 3244 7866 3284 7951
rect 3340 7841 3380 8128
rect 3532 8168 3572 9472
rect 3724 9344 3764 9353
rect 3724 8681 3764 9304
rect 3723 8672 3765 8681
rect 3723 8632 3724 8672
rect 3764 8632 3765 8672
rect 3723 8623 3765 8632
rect 4204 8672 4244 10975
rect 4492 10445 4532 10975
rect 4588 10940 4628 10949
rect 4876 10940 4916 12496
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 4971 12487 5013 12496
rect 4972 12402 5012 12487
rect 5164 11024 5204 13336
rect 5260 13327 5300 13336
rect 6892 13376 6932 13385
rect 5260 12536 5300 12545
rect 5452 12536 5492 12545
rect 6124 12536 6164 12545
rect 5300 12496 5452 12536
rect 5260 12487 5300 12496
rect 5452 12487 5492 12496
rect 5740 12496 6124 12536
rect 5259 12284 5301 12293
rect 5259 12244 5260 12284
rect 5300 12244 5301 12284
rect 5259 12235 5301 12244
rect 5260 12150 5300 12235
rect 5740 11948 5780 12496
rect 6124 12487 6164 12496
rect 5740 11899 5780 11908
rect 6796 12368 6836 12377
rect 6315 11696 6357 11705
rect 6315 11656 6316 11696
rect 6356 11656 6357 11696
rect 6315 11647 6357 11656
rect 6700 11696 6740 11705
rect 6796 11696 6836 12328
rect 6740 11656 6836 11696
rect 6700 11647 6740 11656
rect 6316 11562 6356 11647
rect 6892 11033 6932 13336
rect 11212 13376 11252 13385
rect 8812 13217 8852 13302
rect 7084 13208 7124 13217
rect 7084 12881 7124 13168
rect 7180 13208 7220 13217
rect 7083 12872 7125 12881
rect 7083 12832 7084 12872
rect 7124 12832 7125 12872
rect 7083 12823 7125 12832
rect 7180 12461 7220 13168
rect 7371 13208 7413 13217
rect 8236 13208 8276 13217
rect 7371 13168 7372 13208
rect 7412 13168 7413 13208
rect 7371 13159 7413 13168
rect 7660 13168 8236 13208
rect 7372 13074 7412 13159
rect 7276 13040 7316 13049
rect 7276 12788 7316 13000
rect 7564 13040 7604 13049
rect 7276 12748 7412 12788
rect 7372 12629 7412 12748
rect 7371 12620 7413 12629
rect 7371 12580 7372 12620
rect 7412 12580 7413 12620
rect 7371 12571 7413 12580
rect 7564 12545 7604 13000
rect 7660 12704 7700 13168
rect 8236 13159 8276 13168
rect 8811 13208 8853 13217
rect 8811 13168 8812 13208
rect 8852 13168 8853 13208
rect 8811 13159 8853 13168
rect 8908 13208 8948 13217
rect 8812 13040 8852 13049
rect 7851 12872 7893 12881
rect 7851 12832 7852 12872
rect 7892 12832 7893 12872
rect 7851 12823 7893 12832
rect 8427 12872 8469 12881
rect 8427 12832 8428 12872
rect 8468 12832 8469 12872
rect 8427 12823 8469 12832
rect 7660 12655 7700 12664
rect 7275 12536 7317 12545
rect 7275 12496 7276 12536
rect 7316 12496 7317 12536
rect 7275 12487 7317 12496
rect 7468 12536 7508 12545
rect 7179 12452 7221 12461
rect 7179 12412 7180 12452
rect 7220 12412 7221 12452
rect 7179 12403 7221 12412
rect 7180 11192 7220 12403
rect 7276 12402 7316 12487
rect 7276 12284 7316 12293
rect 7276 11705 7316 12244
rect 7275 11696 7317 11705
rect 7275 11656 7276 11696
rect 7316 11656 7317 11696
rect 7275 11647 7317 11656
rect 7468 11453 7508 12496
rect 7563 12536 7605 12545
rect 7563 12496 7564 12536
rect 7604 12496 7605 12536
rect 7563 12487 7605 12496
rect 7852 12536 7892 12823
rect 8428 12620 8468 12823
rect 8428 12571 8468 12580
rect 7852 12487 7892 12496
rect 7948 12536 7988 12547
rect 7948 12461 7988 12496
rect 8812 12461 8852 13000
rect 8908 12881 8948 13168
rect 9483 13208 9525 13217
rect 9483 13168 9484 13208
rect 9524 13168 9525 13208
rect 9483 13159 9525 13168
rect 10156 13208 10196 13217
rect 9099 13124 9141 13133
rect 9004 13084 9100 13124
rect 9140 13084 9141 13124
rect 8907 12872 8949 12881
rect 8907 12832 8908 12872
rect 8948 12832 8949 12872
rect 8907 12823 8949 12832
rect 7947 12452 7989 12461
rect 7947 12412 7948 12452
rect 7988 12412 7989 12452
rect 7947 12403 7989 12412
rect 8811 12452 8853 12461
rect 8811 12412 8812 12452
rect 8852 12412 8853 12452
rect 8811 12403 8853 12412
rect 8715 11864 8757 11873
rect 8715 11824 8716 11864
rect 8756 11824 8757 11864
rect 8715 11815 8757 11824
rect 8716 11730 8756 11815
rect 7564 11696 7604 11705
rect 9004 11696 9044 13084
rect 9099 13075 9141 13084
rect 9100 12990 9140 13075
rect 9484 13074 9524 13159
rect 9963 12620 10005 12629
rect 9963 12580 9964 12620
rect 10004 12580 10005 12620
rect 9963 12571 10005 12580
rect 9100 12536 9140 12545
rect 9100 11873 9140 12496
rect 9964 12536 10004 12571
rect 9964 12485 10004 12496
rect 9292 12284 9332 12293
rect 9196 12244 9292 12284
rect 9099 11864 9141 11873
rect 9099 11824 9100 11864
rect 9140 11824 9141 11864
rect 9099 11815 9141 11824
rect 9004 11656 9140 11696
rect 7467 11444 7509 11453
rect 7467 11404 7468 11444
rect 7508 11404 7509 11444
rect 7467 11395 7509 11404
rect 7564 11369 7604 11656
rect 9004 11528 9044 11537
rect 8907 11444 8949 11453
rect 8907 11404 8908 11444
rect 8948 11404 8949 11444
rect 8907 11395 8949 11404
rect 7563 11360 7605 11369
rect 7563 11320 7564 11360
rect 7604 11320 7605 11360
rect 7563 11311 7605 11320
rect 8715 11360 8757 11369
rect 8715 11320 8716 11360
rect 8756 11320 8757 11360
rect 8715 11311 8757 11320
rect 7180 11143 7220 11152
rect 7467 11108 7509 11117
rect 7467 11068 7468 11108
rect 7508 11068 7509 11108
rect 7467 11059 7509 11068
rect 5164 10975 5204 10984
rect 6028 11024 6068 11033
rect 4628 10900 4916 10940
rect 4588 10891 4628 10900
rect 4491 10436 4533 10445
rect 4491 10396 4492 10436
rect 4532 10396 4533 10436
rect 4491 10387 4533 10396
rect 5259 10436 5301 10445
rect 5259 10396 5260 10436
rect 5300 10396 5301 10436
rect 5259 10387 5301 10396
rect 4492 10268 4532 10387
rect 5260 10302 5300 10387
rect 4492 10219 4532 10228
rect 6028 10193 6068 10984
rect 6891 11024 6933 11033
rect 6891 10984 6892 11024
rect 6932 10984 6933 11024
rect 6891 10975 6933 10984
rect 7468 10974 7508 11059
rect 7851 11024 7893 11033
rect 7851 10984 7852 11024
rect 7892 10984 7893 11024
rect 7851 10975 7893 10984
rect 8716 11024 8756 11311
rect 8716 10975 8756 10984
rect 7852 10890 7892 10975
rect 6123 10352 6165 10361
rect 6123 10312 6124 10352
rect 6164 10312 6165 10352
rect 6123 10303 6165 10312
rect 6316 10352 6356 10361
rect 6892 10352 6932 10361
rect 4972 10184 5012 10193
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 4204 8623 4244 8632
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4876 8199 4916 8208
rect 3532 8119 3572 8128
rect 4588 8159 4876 8168
rect 4588 8128 4916 8159
rect 4204 8000 4244 8009
rect 4108 7960 4204 8000
rect 4108 7916 4148 7960
rect 4204 7951 4244 7960
rect 4395 8000 4437 8009
rect 4395 7960 4396 8000
rect 4436 7960 4437 8000
rect 4395 7951 4437 7960
rect 4012 7876 4148 7916
rect 1612 7832 1652 7841
rect 1516 7792 1612 7832
rect 1131 7748 1173 7757
rect 1131 7708 1132 7748
rect 1172 7708 1173 7748
rect 1131 7699 1173 7708
rect 1132 7160 1172 7699
rect 1132 7111 1172 7120
rect 1516 7160 1556 7792
rect 1612 7783 1652 7792
rect 3339 7832 3381 7841
rect 3339 7792 3340 7832
rect 3380 7792 3381 7832
rect 3339 7783 3381 7792
rect 2187 7748 2229 7757
rect 2187 7708 2188 7748
rect 2228 7708 2229 7748
rect 2187 7699 2229 7708
rect 2188 7614 2228 7699
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 1516 7111 1556 7120
rect 2380 7160 2420 7169
rect 1420 5816 1460 5825
rect 1324 5776 1420 5816
rect 940 4976 980 4985
rect 940 4397 980 4936
rect 1324 4976 1364 5776
rect 1420 5767 1460 5776
rect 1995 5060 2037 5069
rect 1995 5020 1996 5060
rect 2036 5020 2037 5060
rect 1995 5011 2037 5020
rect 1324 4927 1364 4936
rect 939 4388 981 4397
rect 939 4348 940 4388
rect 980 4348 981 4388
rect 939 4339 981 4348
rect 1611 4388 1653 4397
rect 1611 4348 1612 4388
rect 1652 4348 1653 4388
rect 1611 4339 1653 4348
rect 1612 4254 1652 4339
rect 1707 4136 1749 4145
rect 1707 4096 1708 4136
rect 1748 4096 1749 4136
rect 1707 4087 1749 4096
rect 1708 4002 1748 4087
rect 1996 2624 2036 5011
rect 2380 4985 2420 7120
rect 3532 6992 3572 7001
rect 3532 6749 3572 6952
rect 4012 6749 4052 7876
rect 4203 7832 4245 7841
rect 4203 7792 4204 7832
rect 4244 7792 4245 7832
rect 4203 7783 4245 7792
rect 4396 7832 4436 7951
rect 4396 7783 4436 7792
rect 4108 6992 4148 7001
rect 3531 6740 3573 6749
rect 3531 6700 3532 6740
rect 3572 6700 3573 6740
rect 3531 6691 3573 6700
rect 4011 6740 4053 6749
rect 4011 6700 4012 6740
rect 4052 6700 4053 6740
rect 4011 6691 4053 6700
rect 4108 6497 4148 6952
rect 2667 6488 2709 6497
rect 2667 6448 2668 6488
rect 2708 6448 2709 6488
rect 2667 6439 2709 6448
rect 3052 6488 3092 6497
rect 2668 6354 2708 6439
rect 3052 6320 3092 6448
rect 2956 6280 3092 6320
rect 3916 6488 3956 6497
rect 3916 6320 3956 6448
rect 4107 6488 4149 6497
rect 4107 6448 4108 6488
rect 4148 6448 4149 6488
rect 4107 6439 4149 6448
rect 4204 6320 4244 7783
rect 4588 6992 4628 8128
rect 4972 8084 5012 10144
rect 5932 10184 5972 10193
rect 6027 10184 6069 10193
rect 5972 10144 6028 10184
rect 6068 10144 6069 10184
rect 5932 10135 5972 10144
rect 6027 10135 6069 10144
rect 6028 10050 6068 10135
rect 5548 9640 5972 9680
rect 5260 9512 5300 9521
rect 5452 9512 5492 9521
rect 5548 9512 5588 9640
rect 5300 9472 5396 9512
rect 5260 9463 5300 9472
rect 5356 8924 5396 9472
rect 5492 9472 5588 9512
rect 5644 9512 5684 9521
rect 5452 9463 5492 9472
rect 5452 9344 5492 9353
rect 5644 9344 5684 9472
rect 5492 9304 5684 9344
rect 5452 9295 5492 9304
rect 5548 8924 5588 8933
rect 5356 8884 5548 8924
rect 5548 8875 5588 8884
rect 5644 8672 5684 8681
rect 5548 8632 5644 8672
rect 5356 8504 5396 8513
rect 4876 8044 5012 8084
rect 5068 8464 5356 8504
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4780 8000 4820 8009
rect 4684 7866 4724 7951
rect 4780 7421 4820 7960
rect 4876 7757 4916 8044
rect 5068 8000 5108 8464
rect 5356 8455 5396 8464
rect 5068 7951 5108 7960
rect 5548 7841 5588 8632
rect 5644 8623 5684 8632
rect 5836 8588 5876 8597
rect 5739 8000 5781 8009
rect 5739 7960 5740 8000
rect 5780 7960 5781 8000
rect 5739 7951 5781 7960
rect 5547 7832 5589 7841
rect 5547 7792 5548 7832
rect 5588 7792 5589 7832
rect 5547 7783 5589 7792
rect 4875 7748 4917 7757
rect 4875 7708 4876 7748
rect 4916 7708 4917 7748
rect 4875 7699 4917 7708
rect 4779 7412 4821 7421
rect 4779 7372 4780 7412
rect 4820 7372 4821 7412
rect 4779 7363 4821 7372
rect 4780 7169 4820 7254
rect 4779 7160 4821 7169
rect 4779 7120 4780 7160
rect 4820 7120 4821 7160
rect 4779 7111 4821 7120
rect 4588 6952 4820 6992
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 3916 6280 4052 6320
rect 4204 6280 4532 6320
rect 2956 5816 2996 6280
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 3148 5816 3188 5825
rect 2956 5776 3148 5816
rect 3148 5767 3188 5776
rect 3723 5060 3765 5069
rect 3820 5060 3860 5069
rect 3723 5020 3724 5060
rect 3764 5020 3820 5060
rect 3723 5011 3765 5020
rect 3820 5011 3860 5020
rect 4012 4985 4052 6280
rect 4492 5900 4532 6280
rect 4492 5851 4532 5860
rect 4780 5741 4820 6952
rect 4779 5732 4821 5741
rect 4779 5692 4780 5732
rect 4820 5692 4821 5732
rect 4779 5683 4821 5692
rect 4492 5648 4532 5657
rect 4492 5489 4532 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 4780 5648 4820 5683
rect 4684 5514 4724 5599
rect 4780 5597 4820 5608
rect 4491 5480 4533 5489
rect 4491 5440 4492 5480
rect 4532 5440 4533 5480
rect 4491 5431 4533 5440
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 2187 4976 2229 4985
rect 2187 4936 2188 4976
rect 2228 4936 2229 4976
rect 2187 4927 2229 4936
rect 2379 4976 2421 4985
rect 2379 4936 2380 4976
rect 2420 4936 2421 4976
rect 2379 4927 2421 4936
rect 3436 4976 3476 4985
rect 3916 4976 3956 4985
rect 3476 4936 3572 4976
rect 3436 4927 3476 4936
rect 2188 4842 2228 4927
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 2092 4304 2132 4313
rect 2092 2624 2132 4264
rect 2476 4304 2516 4313
rect 2476 3473 2516 4264
rect 2667 4136 2709 4145
rect 2667 4096 2668 4136
rect 2708 4096 2709 4136
rect 2667 4087 2709 4096
rect 3340 4136 3380 4145
rect 3532 4136 3572 4936
rect 3916 4733 3956 4936
rect 4011 4976 4053 4985
rect 4011 4936 4012 4976
rect 4052 4936 4053 4976
rect 4011 4927 4053 4936
rect 4299 4976 4341 4985
rect 4299 4936 4300 4976
rect 4340 4936 4341 4976
rect 4299 4927 4341 4936
rect 3915 4724 3957 4733
rect 3915 4684 3916 4724
rect 3956 4684 3957 4724
rect 3915 4675 3957 4684
rect 3380 4096 3572 4136
rect 3628 4304 3668 4313
rect 3340 4087 3380 4096
rect 2668 4002 2708 4087
rect 2667 3548 2709 3557
rect 2667 3508 2668 3548
rect 2708 3508 2709 3548
rect 2667 3499 2709 3508
rect 2475 3464 2517 3473
rect 2475 3424 2476 3464
rect 2516 3424 2517 3464
rect 2475 3415 2517 3424
rect 2668 3414 2708 3499
rect 3051 3464 3093 3473
rect 3051 3424 3052 3464
rect 3092 3424 3093 3464
rect 3051 3415 3093 3424
rect 3052 3330 3092 3415
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 2380 2624 2420 2633
rect 2092 2584 2380 2624
rect 1996 2575 2036 2584
rect 2380 2575 2420 2584
rect 3244 2624 3284 2635
rect 3244 2549 3284 2584
rect 3243 2540 3285 2549
rect 3243 2500 3244 2540
rect 3284 2500 3285 2540
rect 3243 2491 3285 2500
rect 3148 1952 3188 1961
rect 2956 1912 3148 1952
rect 2956 1289 2996 1912
rect 3148 1903 3188 1912
rect 3532 1952 3572 1961
rect 3628 1952 3668 4264
rect 4012 4136 4052 4927
rect 4300 4145 4340 4927
rect 4491 4724 4533 4733
rect 4491 4684 4492 4724
rect 4532 4684 4533 4724
rect 4491 4675 4533 4684
rect 4492 4590 4532 4675
rect 3916 3464 3956 3473
rect 4012 3464 4052 4096
rect 4299 4136 4341 4145
rect 4299 4096 4300 4136
rect 4340 4096 4341 4136
rect 4299 4087 4341 4096
rect 4876 4136 4916 7699
rect 4971 7412 5013 7421
rect 4971 7372 4972 7412
rect 5012 7372 5013 7412
rect 4971 7363 5013 7372
rect 4972 7278 5012 7363
rect 5451 7160 5493 7169
rect 5451 7120 5452 7160
rect 5492 7120 5493 7160
rect 5451 7111 5493 7120
rect 4972 6992 5012 7001
rect 4972 5900 5012 6952
rect 5068 6329 5108 6414
rect 5163 6404 5205 6413
rect 5163 6364 5164 6404
rect 5204 6364 5205 6404
rect 5163 6355 5205 6364
rect 5067 6320 5109 6329
rect 5067 6280 5068 6320
rect 5108 6280 5109 6320
rect 5067 6271 5109 6280
rect 5164 5900 5204 6355
rect 4972 5860 5108 5900
rect 4971 5732 5013 5741
rect 4971 5692 4972 5732
rect 5012 5692 5013 5732
rect 4971 5683 5013 5692
rect 4972 5648 5012 5683
rect 5068 5657 5108 5860
rect 5164 5851 5204 5860
rect 4972 5597 5012 5608
rect 5067 5648 5109 5657
rect 5067 5608 5068 5648
rect 5108 5608 5109 5648
rect 5067 5599 5109 5608
rect 5164 5648 5204 5657
rect 5164 5153 5204 5608
rect 5452 5564 5492 7111
rect 5548 6992 5588 7783
rect 5740 7748 5780 7951
rect 5740 7244 5780 7708
rect 5836 7412 5876 8548
rect 5932 8168 5972 9640
rect 6028 9512 6068 9521
rect 6124 9512 6164 10303
rect 6068 9472 6164 9512
rect 6028 9463 6068 9472
rect 6316 8840 6356 10312
rect 6796 10312 6892 10352
rect 6796 9344 6836 10312
rect 6892 10303 6932 10312
rect 7275 10352 7317 10361
rect 7275 10312 7276 10352
rect 7316 10312 7317 10352
rect 7275 10303 7317 10312
rect 7276 10218 7316 10303
rect 6891 10184 6933 10193
rect 6891 10144 6892 10184
rect 6932 10144 6933 10184
rect 8908 10184 8948 11395
rect 9004 11117 9044 11488
rect 9003 11108 9045 11117
rect 9003 11068 9004 11108
rect 9044 11068 9045 11108
rect 9003 11059 9045 11068
rect 9003 10184 9045 10193
rect 8908 10144 9004 10184
rect 9044 10144 9045 10184
rect 6891 10135 6933 10144
rect 9003 10135 9045 10144
rect 6892 9512 6932 10135
rect 8139 10100 8181 10109
rect 8139 10060 8140 10100
rect 8180 10060 8181 10100
rect 8139 10051 8181 10060
rect 8140 9512 8180 10051
rect 9004 10050 9044 10135
rect 9100 10016 9140 11656
rect 9196 10184 9236 12244
rect 9292 12235 9332 12244
rect 10059 11864 10101 11873
rect 10059 11824 10060 11864
rect 10100 11824 10101 11864
rect 10059 11815 10101 11824
rect 9676 11696 9716 11705
rect 9292 11656 9676 11696
rect 9292 10352 9332 11656
rect 9676 11647 9716 11656
rect 9963 11696 10005 11705
rect 9963 11656 9964 11696
rect 10004 11656 10005 11696
rect 9963 11647 10005 11656
rect 10060 11696 10100 11815
rect 10060 11647 10100 11656
rect 10156 11696 10196 13168
rect 10348 13208 10388 13219
rect 10348 13133 10388 13168
rect 10540 13208 10580 13217
rect 10347 13124 10389 13133
rect 10347 13084 10348 13124
rect 10388 13084 10389 13124
rect 10347 13075 10389 13084
rect 10540 13049 10580 13168
rect 10924 13208 10964 13219
rect 10924 13133 10964 13168
rect 10923 13124 10965 13133
rect 10923 13084 10924 13124
rect 10964 13084 10965 13124
rect 10923 13075 10965 13084
rect 10444 13040 10484 13049
rect 10444 12629 10484 13000
rect 10539 13040 10581 13049
rect 10732 13040 10772 13049
rect 10539 13000 10540 13040
rect 10580 13000 10581 13040
rect 10539 12991 10581 13000
rect 10636 13000 10732 13040
rect 10443 12620 10485 12629
rect 10443 12580 10444 12620
rect 10484 12580 10485 12620
rect 10443 12571 10485 12580
rect 9867 11444 9909 11453
rect 9867 11404 9868 11444
rect 9908 11404 9909 11444
rect 9867 11395 9909 11404
rect 9868 11192 9908 11395
rect 9964 11369 10004 11647
rect 10156 11453 10196 11656
rect 10348 12536 10388 12545
rect 10155 11444 10197 11453
rect 10155 11404 10156 11444
rect 10196 11404 10197 11444
rect 10155 11395 10197 11404
rect 9963 11360 10005 11369
rect 9963 11320 9964 11360
rect 10004 11320 10005 11360
rect 9963 11311 10005 11320
rect 9868 11143 9908 11152
rect 9579 10772 9621 10781
rect 9579 10732 9580 10772
rect 9620 10732 9621 10772
rect 9579 10723 9621 10732
rect 9292 10303 9332 10312
rect 9196 10135 9236 10144
rect 9292 10184 9332 10193
rect 9292 10016 9332 10144
rect 9483 10184 9525 10193
rect 9580 10184 9620 10723
rect 9867 10352 9909 10361
rect 9867 10312 9868 10352
rect 9908 10312 9909 10352
rect 9867 10303 9909 10312
rect 9772 10193 9812 10278
rect 9483 10144 9484 10184
rect 9524 10144 9580 10184
rect 9483 10135 9525 10144
rect 9580 10135 9620 10144
rect 9771 10184 9813 10193
rect 9771 10144 9772 10184
rect 9812 10144 9813 10184
rect 9771 10135 9813 10144
rect 9868 10184 9908 10303
rect 9868 10135 9908 10144
rect 9675 10100 9717 10109
rect 9675 10060 9676 10100
rect 9716 10060 9717 10100
rect 9675 10051 9717 10060
rect 9100 9976 9332 10016
rect 9483 10016 9525 10025
rect 9483 9976 9484 10016
rect 9524 9976 9525 10016
rect 9483 9967 9525 9976
rect 6932 9472 7124 9512
rect 6892 9463 6932 9472
rect 6796 9304 6932 9344
rect 6220 8800 6356 8840
rect 6220 8672 6260 8800
rect 6220 8623 6260 8632
rect 5932 8119 5972 8128
rect 5836 7363 5876 7372
rect 6604 8000 6644 8009
rect 6604 7253 6644 7960
rect 6795 7832 6837 7841
rect 6795 7792 6796 7832
rect 6836 7792 6837 7832
rect 6795 7783 6837 7792
rect 6796 7698 6836 7783
rect 6027 7244 6069 7253
rect 5740 7204 5876 7244
rect 5644 7160 5684 7169
rect 5684 7120 5780 7160
rect 5644 7111 5684 7120
rect 5548 6952 5684 6992
rect 5547 6488 5589 6497
rect 5547 6448 5548 6488
rect 5588 6448 5589 6488
rect 5547 6439 5589 6448
rect 5644 6488 5684 6952
rect 5644 6439 5684 6448
rect 5548 6354 5588 6439
rect 5740 6329 5780 7120
rect 5739 6320 5781 6329
rect 5739 6280 5740 6320
rect 5780 6280 5781 6320
rect 5739 6271 5781 6280
rect 5643 5732 5685 5741
rect 5643 5692 5644 5732
rect 5684 5692 5685 5732
rect 5643 5683 5685 5692
rect 5644 5648 5684 5683
rect 5644 5597 5684 5608
rect 5452 5515 5492 5524
rect 5836 5489 5876 7204
rect 6027 7204 6028 7244
rect 6068 7204 6069 7244
rect 6027 7195 6069 7204
rect 6603 7244 6645 7253
rect 6603 7204 6604 7244
rect 6644 7204 6645 7244
rect 6603 7195 6645 7204
rect 5931 7160 5973 7169
rect 5931 7120 5932 7160
rect 5972 7120 5973 7160
rect 5931 7111 5973 7120
rect 5932 6656 5972 7111
rect 5932 6607 5972 6616
rect 6028 6497 6068 7195
rect 6507 7160 6549 7169
rect 6507 7120 6508 7160
rect 6548 7120 6549 7160
rect 6507 7111 6549 7120
rect 6508 7026 6548 7111
rect 6700 6992 6740 7001
rect 6604 6952 6700 6992
rect 6604 6740 6644 6952
rect 6700 6943 6740 6952
rect 6412 6700 6644 6740
rect 6027 6488 6069 6497
rect 6027 6448 6028 6488
rect 6068 6448 6069 6488
rect 6027 6439 6069 6448
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 6412 6488 6452 6700
rect 6507 6572 6549 6581
rect 6507 6532 6508 6572
rect 6548 6532 6549 6572
rect 6507 6523 6549 6532
rect 6412 6439 6452 6448
rect 6028 5900 6068 6439
rect 6220 6354 6260 6439
rect 6315 6320 6357 6329
rect 6508 6320 6548 6523
rect 6796 6488 6836 6497
rect 6892 6488 6932 9304
rect 7084 8672 7124 9472
rect 8140 9463 8180 9472
rect 8524 9512 8564 9521
rect 8524 8849 8564 9472
rect 8908 9512 8948 9521
rect 8948 9472 9044 9512
rect 8908 9463 8948 9472
rect 8523 8840 8565 8849
rect 8523 8800 8524 8840
rect 8564 8800 8565 8840
rect 8523 8791 8565 8800
rect 9004 8840 9044 9472
rect 9004 8791 9044 8800
rect 9387 8840 9429 8849
rect 9387 8800 9388 8840
rect 9428 8800 9429 8840
rect 9387 8791 9429 8800
rect 9388 8706 9428 8791
rect 7084 8623 7124 8632
rect 9484 8672 9524 9967
rect 9676 9966 9716 10051
rect 9964 10016 10004 11311
rect 10060 11024 10100 11033
rect 10060 10277 10100 10984
rect 10348 10520 10388 12496
rect 10444 11528 10484 11537
rect 10444 11369 10484 11488
rect 10443 11360 10485 11369
rect 10443 11320 10444 11360
rect 10484 11320 10485 11360
rect 10443 11311 10485 11320
rect 10539 10772 10581 10781
rect 10539 10732 10540 10772
rect 10580 10732 10581 10772
rect 10539 10723 10581 10732
rect 10348 10480 10484 10520
rect 10059 10268 10101 10277
rect 10059 10228 10060 10268
rect 10100 10228 10101 10268
rect 10059 10219 10101 10228
rect 10251 10268 10293 10277
rect 10251 10228 10252 10268
rect 10292 10228 10293 10268
rect 10251 10219 10293 10228
rect 10156 10184 10196 10195
rect 10156 10109 10196 10144
rect 10252 10184 10292 10219
rect 10155 10100 10197 10109
rect 10155 10060 10156 10100
rect 10196 10060 10197 10100
rect 10155 10051 10197 10060
rect 9772 9976 10004 10016
rect 10059 10016 10101 10025
rect 10059 9976 10060 10016
rect 10100 9976 10101 10016
rect 9772 9512 9812 9976
rect 10059 9967 10101 9976
rect 10060 9882 10100 9967
rect 9772 9463 9812 9472
rect 9484 8623 9524 8632
rect 10252 8672 10292 10144
rect 10347 10184 10389 10193
rect 10347 10144 10348 10184
rect 10388 10144 10389 10184
rect 10347 10135 10389 10144
rect 10348 10050 10388 10135
rect 10347 9428 10389 9437
rect 10347 9388 10348 9428
rect 10388 9388 10389 9428
rect 10347 9379 10389 9388
rect 10252 8623 10292 8632
rect 10348 8672 10388 9379
rect 10444 8840 10484 10480
rect 10444 8791 10484 8800
rect 10348 8623 10388 8632
rect 10540 8672 10580 10723
rect 10636 10277 10676 13000
rect 10732 12991 10772 13000
rect 11019 13040 11061 13049
rect 11019 13000 11020 13040
rect 11060 13000 11061 13040
rect 11019 12991 11061 13000
rect 11020 12906 11060 12991
rect 10732 12536 10772 12545
rect 11212 12536 11252 13336
rect 12364 13208 12404 13217
rect 11691 13040 11733 13049
rect 11691 13000 11692 13040
rect 11732 13000 11733 13040
rect 11691 12991 11733 13000
rect 11692 12906 11732 12991
rect 11499 12620 11541 12629
rect 11499 12580 11500 12620
rect 11540 12580 11541 12620
rect 11499 12571 11541 12580
rect 10772 12496 11252 12536
rect 10732 12487 10772 12496
rect 10828 11696 10868 11705
rect 10731 10772 10773 10781
rect 10731 10732 10732 10772
rect 10772 10732 10773 10772
rect 10731 10723 10773 10732
rect 10732 10638 10772 10723
rect 10635 10268 10677 10277
rect 10635 10228 10636 10268
rect 10676 10228 10677 10268
rect 10635 10219 10677 10228
rect 10731 10184 10773 10193
rect 10731 10144 10732 10184
rect 10772 10144 10773 10184
rect 10731 10135 10773 10144
rect 10732 10050 10772 10135
rect 10540 8623 10580 8632
rect 8236 8504 8276 8513
rect 8236 8009 8276 8464
rect 9100 8084 9140 8093
rect 7467 8000 7509 8009
rect 7467 7960 7468 8000
rect 7508 7960 7509 8000
rect 7467 7951 7509 7960
rect 7756 8000 7796 8009
rect 7468 7866 7508 7951
rect 7372 7160 7412 7169
rect 6836 6448 6932 6488
rect 7275 6488 7317 6497
rect 7275 6448 7276 6488
rect 7316 6448 7317 6488
rect 6796 6439 6836 6448
rect 7275 6439 7317 6448
rect 6315 6280 6316 6320
rect 6356 6280 6357 6320
rect 6315 6271 6357 6280
rect 6412 6280 6548 6320
rect 6123 6236 6165 6245
rect 6123 6196 6124 6236
rect 6164 6196 6165 6236
rect 6123 6187 6165 6196
rect 6124 6102 6164 6187
rect 6220 5900 6260 5909
rect 6028 5860 6220 5900
rect 6220 5851 6260 5860
rect 5931 5648 5973 5657
rect 5931 5608 5932 5648
rect 5972 5608 5973 5648
rect 5931 5599 5973 5608
rect 5932 5514 5972 5599
rect 6316 5564 6356 6271
rect 6412 5648 6452 6280
rect 6795 6236 6837 6245
rect 6795 6196 6796 6236
rect 6836 6196 6837 6236
rect 6795 6187 6837 6196
rect 6508 5741 6548 5772
rect 6507 5732 6549 5741
rect 6507 5692 6508 5732
rect 6548 5692 6549 5732
rect 6507 5683 6549 5692
rect 6412 5599 6452 5608
rect 6508 5648 6548 5683
rect 6316 5515 6356 5524
rect 6508 5489 6548 5608
rect 6603 5648 6645 5657
rect 6603 5608 6604 5648
rect 6644 5608 6645 5648
rect 6603 5599 6645 5608
rect 6796 5648 6836 6187
rect 7276 5909 7316 6439
rect 7372 6413 7412 7120
rect 7563 7160 7605 7169
rect 7563 7120 7564 7160
rect 7604 7120 7605 7160
rect 7563 7111 7605 7120
rect 7467 7076 7509 7085
rect 7467 7036 7468 7076
rect 7508 7036 7509 7076
rect 7467 7027 7509 7036
rect 7371 6404 7413 6413
rect 7371 6364 7372 6404
rect 7412 6364 7413 6404
rect 7371 6355 7413 6364
rect 7275 5900 7317 5909
rect 7275 5860 7276 5900
rect 7316 5860 7412 5900
rect 7275 5851 7317 5860
rect 7084 5648 7124 5657
rect 7276 5648 7316 5657
rect 6836 5608 6932 5648
rect 6796 5599 6836 5608
rect 5835 5480 5877 5489
rect 5835 5440 5836 5480
rect 5876 5440 5877 5480
rect 5835 5431 5877 5440
rect 6219 5480 6261 5489
rect 6219 5440 6220 5480
rect 6260 5440 6261 5480
rect 6219 5431 6261 5440
rect 6507 5480 6549 5489
rect 6507 5440 6508 5480
rect 6548 5440 6549 5480
rect 6507 5431 6549 5440
rect 6220 5346 6260 5431
rect 5163 5144 5205 5153
rect 5163 5104 5164 5144
rect 5204 5104 5205 5144
rect 5163 5095 5205 5104
rect 5356 5148 5396 5157
rect 5164 4976 5204 4985
rect 4971 4724 5013 4733
rect 4971 4684 4972 4724
rect 5012 4684 5013 4724
rect 4971 4675 5013 4684
rect 4876 4087 4916 4096
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 4875 3800 4917 3809
rect 4875 3760 4876 3800
rect 4916 3760 4917 3800
rect 4875 3751 4917 3760
rect 4779 3716 4821 3725
rect 4779 3676 4780 3716
rect 4820 3676 4821 3716
rect 4779 3667 4821 3676
rect 3956 3424 4052 3464
rect 3819 2540 3861 2549
rect 3916 2540 3956 3424
rect 4395 3380 4437 3389
rect 4395 3340 4396 3380
rect 4436 3340 4437 3380
rect 4395 3331 4437 3340
rect 4396 2876 4436 3331
rect 4396 2827 4436 2836
rect 4780 2876 4820 3667
rect 4876 3389 4916 3751
rect 4875 3380 4917 3389
rect 4875 3340 4876 3380
rect 4916 3340 4917 3380
rect 4875 3331 4917 3340
rect 4875 3128 4917 3137
rect 4875 3088 4876 3128
rect 4916 3088 4917 3128
rect 4875 3079 4917 3088
rect 4780 2801 4820 2836
rect 4779 2792 4821 2801
rect 4779 2752 4780 2792
rect 4820 2752 4821 2792
rect 4779 2743 4821 2752
rect 4780 2624 4820 2633
rect 4876 2624 4916 3079
rect 4820 2584 4916 2624
rect 4972 2624 5012 4675
rect 5164 3809 5204 4936
rect 5356 4733 5396 5108
rect 6028 5144 6068 5153
rect 6604 5144 6644 5599
rect 6068 5104 6260 5144
rect 6028 5095 6068 5104
rect 5451 4976 5493 4985
rect 5451 4936 5452 4976
rect 5492 4936 5493 4976
rect 5451 4927 5493 4936
rect 5548 4976 5588 4985
rect 5452 4842 5492 4927
rect 5355 4724 5397 4733
rect 5355 4684 5356 4724
rect 5396 4684 5397 4724
rect 5355 4675 5397 4684
rect 5548 4304 5588 4936
rect 6124 4976 6164 4985
rect 5836 4808 5876 4817
rect 6124 4808 6164 4936
rect 5876 4768 6164 4808
rect 5836 4759 5876 4768
rect 5452 4264 5588 4304
rect 5452 4052 5492 4264
rect 5547 4136 5589 4145
rect 6124 4136 6164 4145
rect 5547 4096 5548 4136
rect 5588 4096 5589 4136
rect 5547 4087 5589 4096
rect 5644 4096 6124 4136
rect 5260 4012 5452 4052
rect 5163 3800 5205 3809
rect 5163 3760 5164 3800
rect 5204 3760 5205 3800
rect 5163 3751 5205 3760
rect 5067 3632 5109 3641
rect 5067 3592 5068 3632
rect 5108 3592 5109 3632
rect 5067 3583 5109 3592
rect 5068 3498 5108 3583
rect 5260 3548 5300 4012
rect 5452 4003 5492 4012
rect 5548 3632 5588 4087
rect 5644 3641 5684 4096
rect 6124 4087 6164 4096
rect 6220 3725 6260 5104
rect 6604 5095 6644 5104
rect 6699 5060 6741 5069
rect 6699 5020 6700 5060
rect 6740 5020 6741 5060
rect 6699 5011 6741 5020
rect 6507 4976 6549 4985
rect 6507 4936 6508 4976
rect 6548 4936 6549 4976
rect 6507 4927 6549 4936
rect 6700 4976 6740 5011
rect 6508 4842 6548 4927
rect 6700 4925 6740 4936
rect 6796 4976 6836 4987
rect 6892 4985 6932 5608
rect 7124 5608 7220 5648
rect 7084 5599 7124 5608
rect 7083 5480 7125 5489
rect 7083 5440 7084 5480
rect 7124 5440 7125 5480
rect 7083 5431 7125 5440
rect 7084 5346 7124 5431
rect 6987 5144 7029 5153
rect 6987 5104 6988 5144
rect 7028 5104 7029 5144
rect 6987 5095 7029 5104
rect 6988 5060 7028 5095
rect 7180 5069 7220 5608
rect 6988 5009 7028 5020
rect 7179 5060 7221 5069
rect 7179 5020 7180 5060
rect 7220 5020 7221 5060
rect 7179 5011 7221 5020
rect 6796 4901 6836 4936
rect 6891 4976 6933 4985
rect 6891 4936 6892 4976
rect 6932 4936 6933 4976
rect 6891 4927 6933 4936
rect 6795 4892 6837 4901
rect 6795 4852 6796 4892
rect 6836 4852 6837 4892
rect 6795 4843 6837 4852
rect 6316 4724 6356 4733
rect 6219 3716 6261 3725
rect 6219 3676 6220 3716
rect 6260 3676 6261 3716
rect 6219 3667 6261 3676
rect 6316 3641 6356 4684
rect 6508 4136 6548 4145
rect 7180 4136 7220 5011
rect 7276 4901 7316 5608
rect 7275 4892 7317 4901
rect 7275 4852 7276 4892
rect 7316 4852 7317 4892
rect 7275 4843 7317 4852
rect 7275 4136 7317 4145
rect 6548 4096 6644 4136
rect 7180 4096 7276 4136
rect 7316 4096 7317 4136
rect 6508 4087 6548 4096
rect 6412 3968 6452 3977
rect 6452 3928 6548 3968
rect 6412 3919 6452 3928
rect 5452 3592 5588 3632
rect 5643 3632 5685 3641
rect 5643 3592 5644 3632
rect 5684 3592 5685 3632
rect 5452 3548 5492 3592
rect 5643 3583 5685 3592
rect 6315 3632 6357 3641
rect 6315 3592 6316 3632
rect 6356 3592 6357 3632
rect 6315 3583 6357 3592
rect 5164 3508 5300 3548
rect 5356 3508 5492 3548
rect 4780 2575 4820 2584
rect 4972 2575 5012 2584
rect 5068 2624 5108 2633
rect 5164 2624 5204 3508
rect 5356 3464 5396 3508
rect 5548 3464 5588 3473
rect 5356 3137 5396 3424
rect 5452 3422 5492 3431
rect 5451 3382 5452 3389
rect 5492 3382 5493 3389
rect 5451 3380 5493 3382
rect 5451 3340 5452 3380
rect 5492 3340 5493 3380
rect 5451 3331 5493 3340
rect 5452 3287 5492 3331
rect 5355 3128 5397 3137
rect 5355 3088 5356 3128
rect 5396 3088 5397 3128
rect 5355 3079 5397 3088
rect 5548 2960 5588 3424
rect 5644 3464 5684 3583
rect 5644 3415 5684 3424
rect 6124 3464 6164 3492
rect 6508 3473 6548 3928
rect 6604 3800 6644 4096
rect 7275 4087 7317 4096
rect 7372 4136 7412 5860
rect 7468 5648 7508 7027
rect 7468 5599 7508 5608
rect 7564 4388 7604 7111
rect 7660 6488 7700 6499
rect 7660 6413 7700 6448
rect 7659 6404 7701 6413
rect 7659 6364 7660 6404
rect 7700 6364 7701 6404
rect 7659 6355 7701 6364
rect 7659 5480 7701 5489
rect 7659 5440 7660 5480
rect 7700 5440 7701 5480
rect 7659 5431 7701 5440
rect 7660 4976 7700 5431
rect 7660 4927 7700 4936
rect 7564 4339 7604 4348
rect 7372 4087 7412 4096
rect 6700 3968 6740 3977
rect 7276 3968 7316 4087
rect 7467 3968 7509 3977
rect 6740 3928 7028 3968
rect 7276 3928 7412 3968
rect 6700 3919 6740 3928
rect 6604 3760 6740 3800
rect 6604 3548 6644 3557
rect 6315 3464 6357 3473
rect 6164 3424 6316 3464
rect 6356 3424 6357 3464
rect 6124 3415 6164 3424
rect 5835 3296 5877 3305
rect 5835 3256 5836 3296
rect 5876 3256 5877 3296
rect 5835 3247 5877 3256
rect 5836 3162 5876 3247
rect 5260 2920 5588 2960
rect 5260 2876 5300 2920
rect 5260 2827 5300 2836
rect 5355 2792 5397 2801
rect 5355 2752 5356 2792
rect 5396 2752 5397 2792
rect 5355 2743 5397 2752
rect 5108 2584 5204 2624
rect 5068 2575 5108 2584
rect 3819 2500 3820 2540
rect 3860 2500 3956 2540
rect 3819 2491 3861 2500
rect 3820 1961 3860 2491
rect 5260 2456 5300 2465
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 3572 1912 3668 1952
rect 3819 1952 3861 1961
rect 3819 1912 3820 1952
rect 3860 1912 3861 1952
rect 3532 1903 3572 1912
rect 3819 1903 3861 1912
rect 4395 1952 4437 1961
rect 4395 1912 4396 1952
rect 4436 1912 4437 1952
rect 4395 1903 4437 1912
rect 4396 1818 4436 1903
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 2955 1280 2997 1289
rect 2955 1240 2956 1280
rect 2996 1240 2997 1280
rect 2955 1231 2997 1240
rect 4107 1280 4149 1289
rect 4107 1240 4108 1280
rect 4148 1240 4149 1280
rect 4107 1231 4149 1240
rect 4108 1146 4148 1231
rect 4972 1196 5012 1205
rect 4780 1156 4972 1196
rect 4780 1112 4820 1156
rect 4972 1147 5012 1156
rect 4780 1063 4820 1072
rect 5260 1112 5300 2416
rect 5260 1063 5300 1072
rect 5356 1112 5396 2743
rect 5932 2624 5972 2633
rect 6124 2624 6164 2633
rect 5548 2584 5932 2624
rect 5548 2120 5588 2584
rect 5932 2575 5972 2584
rect 6028 2584 6124 2624
rect 5548 2071 5588 2080
rect 5932 2120 5972 2129
rect 6028 2120 6068 2584
rect 6124 2575 6164 2584
rect 6220 2549 6260 3424
rect 6315 3415 6357 3424
rect 6412 3464 6452 3473
rect 6316 3396 6356 3415
rect 6412 3305 6452 3424
rect 6507 3464 6549 3473
rect 6507 3424 6508 3464
rect 6548 3424 6549 3464
rect 6507 3415 6549 3424
rect 6411 3296 6453 3305
rect 6411 3256 6412 3296
rect 6452 3256 6453 3296
rect 6411 3247 6453 3256
rect 6604 2633 6644 3508
rect 6700 3305 6740 3760
rect 6988 3690 7028 3928
rect 6988 3473 7028 3650
rect 7083 3548 7125 3557
rect 7083 3508 7084 3548
rect 7124 3508 7125 3548
rect 7083 3499 7125 3508
rect 7275 3548 7317 3557
rect 7275 3508 7276 3548
rect 7316 3508 7317 3548
rect 7275 3499 7317 3508
rect 6987 3464 7029 3473
rect 6987 3424 6988 3464
rect 7028 3424 7029 3464
rect 6987 3415 7029 3424
rect 7084 3464 7124 3499
rect 7084 3413 7124 3424
rect 7180 3464 7220 3475
rect 7180 3389 7220 3424
rect 7179 3380 7221 3389
rect 7179 3340 7180 3380
rect 7220 3340 7221 3380
rect 7179 3331 7221 3340
rect 6699 3296 6741 3305
rect 6699 3256 6700 3296
rect 6740 3256 6741 3296
rect 6699 3247 6741 3256
rect 6987 3296 7029 3305
rect 6987 3256 6988 3296
rect 7028 3256 7029 3296
rect 6987 3247 7029 3256
rect 6603 2624 6645 2633
rect 6603 2584 6604 2624
rect 6644 2584 6645 2624
rect 6603 2575 6645 2584
rect 6988 2624 7028 3247
rect 7180 3128 7220 3331
rect 6988 2575 7028 2584
rect 7084 3088 7220 3128
rect 7084 2624 7124 3088
rect 7084 2575 7124 2584
rect 6219 2540 6261 2549
rect 6219 2500 6220 2540
rect 6260 2500 6261 2540
rect 6219 2491 6261 2500
rect 6795 2540 6837 2549
rect 6795 2500 6796 2540
rect 6836 2500 6837 2540
rect 6795 2491 6837 2500
rect 7179 2540 7221 2549
rect 7179 2500 7180 2540
rect 7220 2500 7221 2540
rect 7179 2491 7221 2500
rect 6796 2406 6836 2491
rect 7180 2406 7220 2491
rect 7276 2456 7316 3499
rect 7276 2407 7316 2416
rect 7372 2456 7412 3928
rect 7467 3928 7468 3968
rect 7508 3928 7509 3968
rect 7467 3919 7509 3928
rect 7468 3296 7508 3919
rect 7756 3893 7796 7960
rect 8235 8000 8277 8009
rect 8235 7960 8236 8000
rect 8276 7960 8277 8000
rect 8235 7951 8277 7960
rect 8715 8000 8757 8009
rect 8715 7960 8716 8000
rect 8756 7960 8757 8000
rect 8715 7951 8757 7960
rect 8139 7916 8181 7925
rect 8139 7876 8140 7916
rect 8180 7876 8181 7916
rect 8139 7867 8181 7876
rect 8043 7748 8085 7757
rect 8043 7708 8044 7748
rect 8084 7708 8085 7748
rect 8043 7699 8085 7708
rect 8044 7614 8084 7699
rect 7852 6992 7892 7001
rect 7852 5060 7892 6952
rect 8140 6320 8180 7867
rect 8716 7866 8756 7951
rect 9100 7244 9140 8044
rect 9196 8000 9236 8011
rect 9196 7925 9236 7960
rect 9580 8000 9620 8009
rect 9195 7916 9237 7925
rect 9195 7876 9196 7916
rect 9236 7876 9237 7916
rect 9195 7867 9237 7876
rect 9580 7337 9620 7960
rect 10156 8000 10196 8011
rect 10828 8009 10868 11656
rect 11403 11024 11445 11033
rect 11403 10984 11404 11024
rect 11444 10984 11445 11024
rect 11500 11024 11540 12571
rect 11596 12536 11636 12545
rect 11596 11696 11636 12496
rect 12267 12368 12309 12377
rect 12267 12328 12268 12368
rect 12308 12328 12309 12368
rect 12267 12319 12309 12328
rect 12075 12284 12117 12293
rect 12075 12244 12076 12284
rect 12116 12244 12117 12284
rect 12075 12235 12117 12244
rect 11691 11696 11733 11705
rect 11596 11656 11692 11696
rect 11732 11656 11733 11696
rect 11691 11647 11733 11656
rect 11692 11562 11732 11647
rect 11884 11612 11924 11621
rect 11691 11360 11733 11369
rect 11691 11320 11692 11360
rect 11732 11320 11733 11360
rect 11691 11311 11733 11320
rect 11596 11024 11636 11033
rect 11500 10984 11596 11024
rect 11403 10975 11445 10984
rect 11596 10975 11636 10984
rect 10924 10772 10964 10781
rect 10924 9437 10964 10732
rect 11307 10772 11349 10781
rect 11307 10732 11308 10772
rect 11348 10732 11349 10772
rect 11307 10723 11349 10732
rect 11019 10184 11061 10193
rect 11019 10144 11020 10184
rect 11060 10144 11061 10184
rect 11019 10135 11061 10144
rect 10923 9428 10965 9437
rect 10923 9388 10924 9428
rect 10964 9388 10965 9428
rect 10923 9379 10965 9388
rect 10924 9260 10964 9269
rect 11020 9260 11060 10135
rect 11211 9596 11253 9605
rect 11211 9556 11212 9596
rect 11252 9556 11253 9596
rect 11211 9547 11253 9556
rect 11212 9462 11252 9547
rect 11308 9512 11348 10723
rect 11404 10193 11444 10975
rect 11403 10184 11445 10193
rect 11403 10144 11404 10184
rect 11444 10144 11445 10184
rect 11692 10184 11732 11311
rect 11787 11024 11829 11033
rect 11787 10984 11788 11024
rect 11828 10984 11829 11024
rect 11787 10975 11829 10984
rect 11788 10890 11828 10975
rect 11884 10781 11924 11572
rect 12076 11024 12116 12235
rect 12268 11696 12308 12319
rect 12364 12293 12404 13168
rect 12939 12368 12981 12377
rect 12939 12328 12940 12368
rect 12980 12328 12981 12368
rect 12939 12319 12981 12328
rect 12363 12284 12405 12293
rect 12363 12244 12364 12284
rect 12404 12244 12405 12284
rect 12363 12235 12405 12244
rect 12747 12284 12789 12293
rect 12747 12244 12748 12284
rect 12788 12244 12789 12284
rect 12747 12235 12789 12244
rect 12748 12150 12788 12235
rect 12940 12234 12980 12319
rect 12268 11647 12308 11656
rect 13131 11696 13173 11705
rect 13131 11656 13132 11696
rect 13172 11656 13173 11696
rect 13131 11647 13173 11656
rect 12268 11108 12308 11117
rect 12076 10975 12116 10984
rect 12172 11068 12268 11108
rect 11883 10772 11925 10781
rect 11883 10732 11884 10772
rect 11924 10732 11925 10772
rect 11883 10723 11925 10732
rect 11788 10184 11828 10193
rect 11692 10144 11788 10184
rect 11403 10135 11445 10144
rect 11788 10135 11828 10144
rect 11884 10184 11924 10193
rect 12172 10184 12212 11068
rect 12268 11059 12308 11068
rect 12364 10352 12404 10361
rect 11924 10144 12212 10184
rect 12268 10312 12364 10352
rect 11884 10135 11924 10144
rect 11404 10050 11444 10135
rect 11596 10016 11636 10025
rect 10964 9220 11060 9260
rect 11308 9260 11348 9472
rect 11404 9512 11444 9523
rect 11404 9437 11444 9472
rect 11499 9512 11541 9521
rect 11499 9472 11500 9512
rect 11540 9472 11541 9512
rect 11499 9463 11541 9472
rect 11403 9428 11445 9437
rect 11403 9388 11404 9428
rect 11444 9388 11445 9428
rect 11403 9379 11445 9388
rect 11500 9378 11540 9463
rect 11596 9437 11636 9976
rect 12171 10016 12213 10025
rect 12171 9976 12172 10016
rect 12212 9976 12213 10016
rect 12171 9967 12213 9976
rect 12172 9596 12212 9967
rect 11788 9512 11828 9521
rect 11595 9428 11637 9437
rect 11595 9388 11596 9428
rect 11636 9388 11637 9428
rect 11595 9379 11637 9388
rect 11788 9260 11828 9472
rect 11883 9512 11925 9521
rect 11883 9472 11884 9512
rect 11924 9472 11925 9512
rect 11883 9463 11925 9472
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 11884 9353 11924 9463
rect 12076 9378 12116 9463
rect 11883 9344 11925 9353
rect 11883 9304 11884 9344
rect 11924 9304 11925 9344
rect 11883 9295 11925 9304
rect 11308 9220 11828 9260
rect 10924 9211 10964 9220
rect 11499 8840 11541 8849
rect 11499 8800 11500 8840
rect 11540 8800 11541 8840
rect 11499 8791 11541 8800
rect 10924 8672 10964 8681
rect 10964 8632 11156 8672
rect 10924 8623 10964 8632
rect 11116 8168 11156 8632
rect 11116 8119 11156 8128
rect 10156 7925 10196 7960
rect 10348 8000 10388 8009
rect 10635 8000 10677 8009
rect 10388 7960 10484 8000
rect 10348 7951 10388 7960
rect 10155 7916 10197 7925
rect 10155 7876 10156 7916
rect 10196 7876 10197 7916
rect 10155 7867 10197 7876
rect 10348 7748 10388 7757
rect 9579 7328 9621 7337
rect 9579 7288 9580 7328
rect 9620 7288 9621 7328
rect 9579 7279 9621 7288
rect 9100 7204 9524 7244
rect 8523 7160 8565 7169
rect 8523 7120 8524 7160
rect 8564 7120 8565 7160
rect 8523 7111 8565 7120
rect 8716 7160 8756 7169
rect 8524 7026 8564 7111
rect 8716 6320 8756 7120
rect 8907 7160 8949 7169
rect 8907 7120 8908 7160
rect 8948 7120 8949 7160
rect 8907 7111 8949 7120
rect 8811 7076 8853 7085
rect 8811 7036 8812 7076
rect 8852 7036 8853 7076
rect 8811 7027 8853 7036
rect 8812 6942 8852 7027
rect 8908 7026 8948 7111
rect 9196 7076 9236 7085
rect 9196 6656 9236 7036
rect 9484 6992 9524 7204
rect 9580 7160 9620 7169
rect 9620 7120 10100 7160
rect 9580 7111 9620 7120
rect 9484 6952 9908 6992
rect 9196 6607 9236 6616
rect 9868 6488 9908 6952
rect 9868 6439 9908 6448
rect 9099 6404 9141 6413
rect 9099 6364 9100 6404
rect 9140 6364 9141 6404
rect 9099 6355 9141 6364
rect 8044 6280 8180 6320
rect 8620 6280 8756 6320
rect 8044 5657 8084 6280
rect 8139 5984 8181 5993
rect 8139 5944 8140 5984
rect 8180 5944 8181 5984
rect 8139 5935 8181 5944
rect 8043 5648 8085 5657
rect 8043 5608 8044 5648
rect 8084 5608 8085 5648
rect 8043 5599 8085 5608
rect 8140 5648 8180 5935
rect 8524 5900 8564 5909
rect 8620 5900 8660 6280
rect 8140 5599 8180 5608
rect 8332 5860 8524 5900
rect 8564 5860 8660 5900
rect 8812 6236 8852 6245
rect 8332 5648 8372 5860
rect 8524 5851 8564 5860
rect 8812 5657 8852 6196
rect 8332 5599 8372 5608
rect 8811 5648 8853 5657
rect 8811 5608 8812 5648
rect 8852 5608 8853 5648
rect 8811 5599 8853 5608
rect 8044 5514 8084 5599
rect 8235 5480 8277 5489
rect 8235 5440 8236 5480
rect 8276 5440 8277 5480
rect 8235 5431 8277 5440
rect 8236 5346 8276 5431
rect 7852 5011 7892 5020
rect 8236 4976 8276 4985
rect 8236 4304 8276 4936
rect 8715 4976 8757 4985
rect 8715 4936 8716 4976
rect 8756 4936 8757 4976
rect 8715 4927 8757 4936
rect 9100 4976 9140 6355
rect 10060 6320 10100 7120
rect 10060 6271 10100 6280
rect 9387 5900 9429 5909
rect 9387 5860 9388 5900
rect 9428 5860 9429 5900
rect 9387 5851 9429 5860
rect 9388 5766 9428 5851
rect 9195 5648 9237 5657
rect 9195 5608 9196 5648
rect 9236 5608 9237 5648
rect 9195 5599 9237 5608
rect 10060 5648 10100 5657
rect 10100 5608 10292 5648
rect 10060 5599 10100 5608
rect 9196 5514 9236 5599
rect 8332 4304 8372 4313
rect 8236 4264 8332 4304
rect 8332 4255 8372 4264
rect 7851 4136 7893 4145
rect 7851 4096 7852 4136
rect 7892 4096 7893 4136
rect 7851 4087 7893 4096
rect 7948 4136 7988 4145
rect 7852 3968 7892 4087
rect 7948 3977 7988 4096
rect 8716 4136 8756 4927
rect 9100 4817 9140 4936
rect 10252 4892 10292 5608
rect 10252 4843 10292 4852
rect 9099 4808 9141 4817
rect 9099 4768 9100 4808
rect 9140 4768 9141 4808
rect 9099 4759 9141 4768
rect 9675 4808 9717 4817
rect 9675 4768 9676 4808
rect 9716 4768 9717 4808
rect 9675 4759 9717 4768
rect 8716 4087 8756 4096
rect 8907 4136 8949 4145
rect 8907 4096 8908 4136
rect 8948 4096 8949 4136
rect 8907 4087 8949 4096
rect 8908 4002 8948 4087
rect 7852 3919 7892 3928
rect 7947 3968 7989 3977
rect 7947 3928 7948 3968
rect 7988 3928 7989 3968
rect 7947 3919 7989 3928
rect 8140 3968 8180 3977
rect 8812 3968 8852 3977
rect 8180 3928 8564 3968
rect 8140 3919 8180 3928
rect 7755 3884 7797 3893
rect 7755 3844 7756 3884
rect 7796 3844 7797 3884
rect 7755 3835 7797 3844
rect 7659 3548 7701 3557
rect 7659 3508 7660 3548
rect 7700 3508 7701 3548
rect 7659 3499 7701 3508
rect 8140 3548 8180 3557
rect 8180 3508 8468 3548
rect 8140 3499 8180 3508
rect 7660 3464 7700 3499
rect 7660 3413 7700 3424
rect 7947 3464 7989 3473
rect 7947 3424 7948 3464
rect 7988 3424 7989 3464
rect 7947 3415 7989 3424
rect 8428 3464 8468 3508
rect 8428 3415 8468 3424
rect 7948 3330 7988 3415
rect 7468 3247 7508 3256
rect 7563 2624 7605 2633
rect 7563 2584 7564 2624
rect 7604 2584 7605 2624
rect 7563 2575 7605 2584
rect 8428 2624 8468 2633
rect 8524 2624 8564 3928
rect 8812 3473 8852 3928
rect 9388 3968 9428 3977
rect 9388 3557 9428 3928
rect 9387 3548 9429 3557
rect 9387 3508 9388 3548
rect 9428 3508 9429 3548
rect 9387 3499 9429 3508
rect 8811 3464 8853 3473
rect 8811 3424 8812 3464
rect 8852 3424 8853 3464
rect 8811 3415 8853 3424
rect 9387 3380 9429 3389
rect 9387 3340 9388 3380
rect 9428 3340 9429 3380
rect 9387 3331 9429 3340
rect 8811 3296 8853 3305
rect 8811 3256 8812 3296
rect 8852 3256 8853 3296
rect 8811 3247 8853 3256
rect 8619 3212 8661 3221
rect 8619 3172 8620 3212
rect 8660 3172 8661 3212
rect 8619 3163 8661 3172
rect 8468 2584 8564 2624
rect 8428 2575 8468 2584
rect 7564 2490 7604 2575
rect 7372 2407 7412 2416
rect 8236 2456 8276 2465
rect 5972 2080 6068 2120
rect 5932 2071 5972 2080
rect 8236 2036 8276 2416
rect 8332 2036 8372 2045
rect 8236 1996 8332 2036
rect 8332 1987 8372 1996
rect 8524 2036 8564 2045
rect 8620 2036 8660 3163
rect 8812 2624 8852 3247
rect 9388 3246 9428 3331
rect 9099 3212 9141 3221
rect 9099 3172 9100 3212
rect 9140 3172 9141 3212
rect 9099 3163 9141 3172
rect 9100 3078 9140 3163
rect 8812 2575 8852 2584
rect 9676 2624 9716 4759
rect 10348 4145 10388 7708
rect 10444 7589 10484 7960
rect 10635 7960 10636 8000
rect 10676 7960 10677 8000
rect 10635 7951 10677 7960
rect 10827 8000 10869 8009
rect 10827 7960 10828 8000
rect 10868 7960 10869 8000
rect 10827 7951 10869 7960
rect 11307 8000 11349 8009
rect 11307 7960 11308 8000
rect 11348 7960 11349 8000
rect 11500 8000 11540 8791
rect 11596 8672 11636 8681
rect 11788 8672 11828 8681
rect 11636 8632 11788 8672
rect 11596 8623 11636 8632
rect 11788 8623 11828 8632
rect 11884 8168 11924 9295
rect 12172 8849 12212 9556
rect 12171 8840 12213 8849
rect 12171 8800 12172 8840
rect 12212 8800 12213 8840
rect 12171 8791 12213 8800
rect 12172 8672 12212 8681
rect 12268 8672 12308 10312
rect 12364 10303 12404 10312
rect 12747 10016 12789 10025
rect 12747 9976 12748 10016
rect 12788 9976 12789 10016
rect 12747 9967 12789 9976
rect 12748 9882 12788 9967
rect 12651 9512 12693 9521
rect 12651 9472 12652 9512
rect 12692 9472 12693 9512
rect 12651 9463 12693 9472
rect 12652 9378 12692 9463
rect 12212 8632 12308 8672
rect 12460 9260 12500 9269
rect 12172 8623 12212 8632
rect 11884 8119 11924 8128
rect 12460 8093 12500 9220
rect 13036 8672 13076 8681
rect 13132 8672 13172 11647
rect 14284 11528 14324 11537
rect 14092 11488 14284 11528
rect 14092 10940 14132 11488
rect 14284 11479 14324 11488
rect 14283 11192 14325 11201
rect 14283 11152 14284 11192
rect 14324 11152 14325 11192
rect 14283 11143 14325 11152
rect 14284 11058 14324 11143
rect 14092 10891 14132 10900
rect 13420 10184 13460 10193
rect 13420 9764 13460 10144
rect 13420 9724 14132 9764
rect 13515 9596 13557 9605
rect 13515 9556 13516 9596
rect 13556 9556 13557 9596
rect 13515 9547 13557 9556
rect 13324 9512 13364 9521
rect 13324 9353 13364 9472
rect 13516 9512 13556 9547
rect 13516 9461 13556 9472
rect 13708 9512 13748 9521
rect 13708 9353 13748 9472
rect 13803 9512 13845 9521
rect 13803 9472 13804 9512
rect 13844 9472 13845 9512
rect 13803 9463 13845 9472
rect 13804 9378 13844 9463
rect 13323 9344 13365 9353
rect 13323 9304 13324 9344
rect 13364 9304 13365 9344
rect 13323 9295 13365 9304
rect 13707 9344 13749 9353
rect 13996 9344 14036 9353
rect 13707 9304 13708 9344
rect 13748 9304 13749 9344
rect 13707 9295 13749 9304
rect 13900 9304 13996 9344
rect 13076 8632 13172 8672
rect 13516 9260 13556 9269
rect 12459 8084 12501 8093
rect 12459 8044 12460 8084
rect 12500 8044 12501 8084
rect 12459 8035 12501 8044
rect 11596 8000 11636 8009
rect 11500 7960 11596 8000
rect 11307 7951 11349 7960
rect 11596 7951 11636 7960
rect 13036 8000 13076 8632
rect 13516 8009 13556 9220
rect 13036 7951 13076 7960
rect 13515 8000 13557 8009
rect 13515 7960 13516 8000
rect 13556 7960 13557 8000
rect 13515 7951 13557 7960
rect 13900 8000 13940 9304
rect 13996 9295 14036 9304
rect 13900 7951 13940 7960
rect 14092 8672 14132 9724
rect 14188 8672 14228 8681
rect 14092 8632 14188 8672
rect 10443 7580 10485 7589
rect 10443 7540 10444 7580
rect 10484 7540 10485 7580
rect 10443 7531 10485 7540
rect 10444 7160 10484 7169
rect 10444 6413 10484 7120
rect 10443 6404 10485 6413
rect 10443 6364 10444 6404
rect 10484 6364 10485 6404
rect 10443 6355 10485 6364
rect 10540 5564 10580 5573
rect 10540 4388 10580 5524
rect 10636 4976 10676 7951
rect 11308 7866 11348 7951
rect 11691 7580 11733 7589
rect 11691 7540 11692 7580
rect 11732 7540 11733 7580
rect 11691 7531 11733 7540
rect 10923 7328 10965 7337
rect 10923 7288 10924 7328
rect 10964 7288 10965 7328
rect 10923 7279 10965 7288
rect 10731 7160 10773 7169
rect 10731 7120 10732 7160
rect 10772 7120 10773 7160
rect 10731 7111 10773 7120
rect 10732 6656 10772 7111
rect 10732 6607 10772 6616
rect 10924 5648 10964 7279
rect 11596 6992 11636 7001
rect 11404 6952 11596 6992
rect 11404 6488 11444 6952
rect 11596 6943 11636 6952
rect 11404 5993 11444 6448
rect 11692 6320 11732 7531
rect 11787 7328 11829 7337
rect 11787 7288 11788 7328
rect 11828 7288 11829 7328
rect 11787 7279 11829 7288
rect 11788 7194 11828 7279
rect 12556 6488 12596 6497
rect 12556 6320 12596 6448
rect 11596 6280 11732 6320
rect 12172 6280 12596 6320
rect 12748 6320 12788 6329
rect 11403 5984 11445 5993
rect 11403 5944 11404 5984
rect 11444 5944 11445 5984
rect 11403 5935 11445 5944
rect 10924 5599 10964 5608
rect 11596 5144 11636 6280
rect 11884 6236 11924 6245
rect 10636 4927 10676 4936
rect 11404 5104 11636 5144
rect 11788 5648 11828 5657
rect 10827 4808 10869 4817
rect 10827 4768 10828 4808
rect 10868 4768 10869 4808
rect 10827 4759 10869 4768
rect 10828 4674 10868 4759
rect 11020 4724 11060 4733
rect 10540 4339 10580 4348
rect 10060 4136 10100 4145
rect 8564 1996 8660 2036
rect 8524 1987 8564 1996
rect 7083 1952 7125 1961
rect 7083 1912 7084 1952
rect 7124 1912 7125 1952
rect 7083 1903 7125 1912
rect 7948 1952 7988 1961
rect 7084 1818 7124 1903
rect 7948 1289 7988 1912
rect 8908 1952 8948 1961
rect 9676 1952 9716 2584
rect 9964 4096 10060 4136
rect 9964 2129 10004 4096
rect 10060 4087 10100 4096
rect 10347 4136 10389 4145
rect 10347 4096 10348 4136
rect 10388 4096 10389 4136
rect 10347 4087 10389 4096
rect 10827 4052 10869 4061
rect 10827 4012 10828 4052
rect 10868 4012 10869 4052
rect 10827 4003 10869 4012
rect 10731 3800 10773 3809
rect 10731 3760 10732 3800
rect 10772 3760 10773 3800
rect 10731 3751 10773 3760
rect 10060 3464 10100 3473
rect 10060 2885 10100 3424
rect 10635 3464 10677 3473
rect 10635 3424 10636 3464
rect 10676 3424 10677 3464
rect 10635 3415 10677 3424
rect 10732 3464 10772 3751
rect 10828 3632 10868 4003
rect 10828 3583 10868 3592
rect 10732 3415 10772 3424
rect 10923 3464 10965 3473
rect 10923 3424 10924 3464
rect 10964 3424 10965 3464
rect 10923 3415 10965 3424
rect 10636 3330 10676 3415
rect 10924 3330 10964 3415
rect 10251 3296 10293 3305
rect 10251 3256 10252 3296
rect 10292 3256 10293 3296
rect 10251 3247 10293 3256
rect 10252 3162 10292 3247
rect 10059 2876 10101 2885
rect 10059 2836 10060 2876
rect 10100 2836 10101 2876
rect 10059 2827 10101 2836
rect 10827 2876 10869 2885
rect 10827 2836 10828 2876
rect 10868 2836 10869 2876
rect 10827 2827 10869 2836
rect 10828 2742 10868 2827
rect 11020 2708 11060 4684
rect 11404 4388 11444 5104
rect 11788 4985 11828 5608
rect 11884 5060 11924 6196
rect 11884 5011 11924 5020
rect 11500 4976 11540 4985
rect 11787 4976 11829 4985
rect 11540 4936 11788 4976
rect 11828 4936 11829 4976
rect 11500 4927 11540 4936
rect 11787 4927 11829 4936
rect 11788 4842 11828 4927
rect 11979 4892 12021 4901
rect 11979 4852 11980 4892
rect 12020 4852 12021 4892
rect 11979 4843 12021 4852
rect 11404 4339 11444 4348
rect 11211 4136 11253 4145
rect 11211 4096 11212 4136
rect 11252 4096 11253 4136
rect 11211 4087 11253 4096
rect 11212 4002 11252 4087
rect 11691 3968 11733 3977
rect 11691 3928 11692 3968
rect 11732 3928 11733 3968
rect 11691 3919 11733 3928
rect 11211 3632 11253 3641
rect 11211 3592 11212 3632
rect 11252 3592 11253 3632
rect 11211 3583 11253 3592
rect 11212 3498 11252 3583
rect 11307 3548 11349 3557
rect 11307 3508 11308 3548
rect 11348 3508 11349 3548
rect 11307 3499 11349 3508
rect 11308 3464 11348 3499
rect 11308 3413 11348 3424
rect 11692 3464 11732 3919
rect 11980 3548 12020 4843
rect 12076 4145 12116 4230
rect 12075 4136 12117 4145
rect 12075 4096 12076 4136
rect 12116 4096 12117 4136
rect 12075 4087 12117 4096
rect 12075 3968 12117 3977
rect 12075 3928 12076 3968
rect 12116 3928 12117 3968
rect 12075 3919 12117 3928
rect 11980 3499 12020 3508
rect 11692 3415 11732 3424
rect 11883 3464 11925 3473
rect 11883 3424 11884 3464
rect 11924 3424 11925 3464
rect 11883 3415 11925 3424
rect 12076 3464 12116 3919
rect 12172 3641 12212 6280
rect 12268 4976 12308 4985
rect 12748 4976 12788 6280
rect 12308 4936 12788 4976
rect 12940 5480 12980 5489
rect 12268 4927 12308 4936
rect 12940 4136 12980 5440
rect 13131 4976 13173 4985
rect 13131 4936 13132 4976
rect 13172 4936 13173 4976
rect 13131 4927 13173 4936
rect 13132 4842 13172 4927
rect 14092 4220 14132 8632
rect 14188 8623 14228 8632
rect 14283 8084 14325 8093
rect 14283 8044 14284 8084
rect 14324 8044 14325 8084
rect 14283 8035 14325 8044
rect 14284 7950 14324 8035
rect 14284 4724 14324 4733
rect 14092 4171 14132 4180
rect 14188 4684 14284 4724
rect 12940 4087 12980 4096
rect 13804 4136 13844 4145
rect 13804 4052 13844 4096
rect 14188 4052 14228 4684
rect 14284 4675 14324 4684
rect 13804 4012 14228 4052
rect 12268 3968 12308 3977
rect 12171 3632 12213 3641
rect 12171 3592 12172 3632
rect 12212 3592 12213 3632
rect 12171 3583 12213 3592
rect 12268 3473 12308 3928
rect 13131 3968 13173 3977
rect 13131 3928 13132 3968
rect 13172 3928 13173 3968
rect 13131 3919 13173 3928
rect 13132 3834 13172 3919
rect 13804 3809 13844 4012
rect 14284 3968 14324 3977
rect 14284 3809 14324 3928
rect 13803 3800 13845 3809
rect 13803 3760 13804 3800
rect 13844 3760 13845 3800
rect 13803 3751 13845 3760
rect 14283 3800 14325 3809
rect 14283 3760 14284 3800
rect 14324 3760 14325 3800
rect 14283 3751 14325 3760
rect 12076 3415 12116 3424
rect 12267 3464 12309 3473
rect 12267 3424 12268 3464
rect 12308 3424 12309 3464
rect 12267 3415 12309 3424
rect 11884 3330 11924 3415
rect 11020 2659 11060 2668
rect 9963 2120 10005 2129
rect 9963 2080 9964 2120
rect 10004 2080 10005 2120
rect 9963 2071 10005 2080
rect 10923 2120 10965 2129
rect 10923 2080 10924 2120
rect 10964 2080 10965 2120
rect 10923 2071 10965 2080
rect 10924 1986 10964 2071
rect 9772 1952 9812 1961
rect 8948 1912 9428 1952
rect 9676 1912 9772 1952
rect 8908 1903 8948 1912
rect 7083 1280 7125 1289
rect 7083 1240 7084 1280
rect 7124 1240 7125 1280
rect 7083 1231 7125 1240
rect 7947 1280 7989 1289
rect 7947 1240 7948 1280
rect 7988 1240 7989 1280
rect 7947 1231 7989 1240
rect 9388 1280 9428 1912
rect 9772 1903 9812 1912
rect 9388 1231 9428 1240
rect 7084 1146 7124 1231
rect 5356 1063 5396 1072
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
<< via2 >>
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 2188 12244 2228 12284
rect 844 11152 884 11192
rect 1900 10984 1940 11024
rect 2764 12244 2804 12284
rect 4108 12496 4148 12536
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3340 11656 3380 11696
rect 4780 12244 4820 12284
rect 4108 11656 4148 11696
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3436 10984 3476 11024
rect 4204 10984 4244 11024
rect 4492 10984 4532 11024
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 3340 8632 3380 8672
rect 3244 7960 3284 8000
rect 3724 8632 3764 8672
rect 4972 12496 5012 12536
rect 5260 12244 5300 12284
rect 6316 11656 6356 11696
rect 7084 12832 7124 12872
rect 7372 13168 7412 13208
rect 7372 12580 7412 12620
rect 8812 13168 8852 13208
rect 7852 12832 7892 12872
rect 8428 12832 8468 12872
rect 7276 12496 7316 12536
rect 7180 12412 7220 12452
rect 7276 11656 7316 11696
rect 7564 12496 7604 12536
rect 9484 13168 9524 13208
rect 9100 13084 9140 13124
rect 8908 12832 8948 12872
rect 7948 12412 7988 12452
rect 8812 12412 8852 12452
rect 8716 11824 8756 11864
rect 9964 12580 10004 12620
rect 9100 11824 9140 11864
rect 7468 11404 7508 11444
rect 8908 11404 8948 11444
rect 7564 11320 7604 11360
rect 8716 11320 8756 11360
rect 7468 11068 7508 11108
rect 4492 10396 4532 10436
rect 5260 10396 5300 10436
rect 6892 10984 6932 11024
rect 7852 10984 7892 11024
rect 6124 10312 6164 10352
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 4396 7960 4436 8000
rect 1132 7708 1172 7748
rect 3340 7792 3380 7832
rect 2188 7708 2228 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 1996 5020 2036 5060
rect 940 4348 980 4388
rect 1612 4348 1652 4388
rect 1708 4096 1748 4136
rect 4204 7792 4244 7832
rect 3532 6700 3572 6740
rect 4012 6700 4052 6740
rect 2668 6448 2708 6488
rect 4108 6448 4148 6488
rect 6028 10144 6068 10184
rect 4684 7960 4724 8000
rect 5740 7960 5780 8000
rect 5548 7792 5588 7832
rect 4876 7708 4916 7748
rect 4780 7372 4820 7412
rect 4780 7120 4820 7160
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 3724 5020 3764 5060
rect 4780 5692 4820 5732
rect 4684 5608 4724 5648
rect 4492 5440 4532 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 2188 4936 2228 4976
rect 2380 4936 2420 4976
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 2668 4096 2708 4136
rect 4012 4936 4052 4976
rect 4300 4936 4340 4976
rect 3916 4684 3956 4724
rect 2668 3508 2708 3548
rect 2476 3424 2516 3464
rect 3052 3424 3092 3464
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 3244 2500 3284 2540
rect 4492 4684 4532 4724
rect 4300 4096 4340 4136
rect 4972 7372 5012 7412
rect 5452 7120 5492 7160
rect 5164 6364 5204 6404
rect 5068 6280 5108 6320
rect 4972 5692 5012 5732
rect 5068 5608 5108 5648
rect 7276 10312 7316 10352
rect 6892 10144 6932 10184
rect 9004 11068 9044 11108
rect 9004 10144 9044 10184
rect 8140 10060 8180 10100
rect 10060 11824 10100 11864
rect 9964 11656 10004 11696
rect 10348 13084 10388 13124
rect 10924 13084 10964 13124
rect 10540 13000 10580 13040
rect 10444 12580 10484 12620
rect 9868 11404 9908 11444
rect 10156 11404 10196 11444
rect 9964 11320 10004 11360
rect 9580 10732 9620 10772
rect 9868 10312 9908 10352
rect 9484 10144 9524 10184
rect 9772 10144 9812 10184
rect 9676 10060 9716 10100
rect 9484 9976 9524 10016
rect 6796 7792 6836 7832
rect 5548 6448 5588 6488
rect 5740 6280 5780 6320
rect 5644 5692 5684 5732
rect 6028 7204 6068 7244
rect 6604 7204 6644 7244
rect 5932 7120 5972 7160
rect 6508 7120 6548 7160
rect 6028 6448 6068 6488
rect 6220 6448 6260 6488
rect 6508 6532 6548 6572
rect 8524 8800 8564 8840
rect 9388 8800 9428 8840
rect 10444 11320 10484 11360
rect 10540 10732 10580 10772
rect 10060 10228 10100 10268
rect 10252 10228 10292 10268
rect 10156 10060 10196 10100
rect 10060 9976 10100 10016
rect 10348 10144 10388 10184
rect 10348 9388 10388 9428
rect 11020 13000 11060 13040
rect 11692 13000 11732 13040
rect 11500 12580 11540 12620
rect 10732 10732 10772 10772
rect 10636 10228 10676 10268
rect 10732 10144 10772 10184
rect 7468 7960 7508 8000
rect 7276 6448 7316 6488
rect 6316 6280 6356 6320
rect 6124 6196 6164 6236
rect 5932 5608 5972 5648
rect 6796 6196 6836 6236
rect 6508 5692 6548 5732
rect 6604 5608 6644 5648
rect 7564 7120 7604 7160
rect 7468 7036 7508 7076
rect 7372 6364 7412 6404
rect 7276 5860 7316 5900
rect 5836 5440 5876 5480
rect 6220 5440 6260 5480
rect 6508 5440 6548 5480
rect 5164 5104 5204 5144
rect 4972 4684 5012 4724
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 4876 3760 4916 3800
rect 4780 3676 4820 3716
rect 4396 3340 4436 3380
rect 4876 3340 4916 3380
rect 4876 3088 4916 3128
rect 4780 2752 4820 2792
rect 5452 4936 5492 4976
rect 5356 4684 5396 4724
rect 5548 4096 5588 4136
rect 5164 3760 5204 3800
rect 5068 3592 5108 3632
rect 6700 5020 6740 5060
rect 6508 4936 6548 4976
rect 7084 5440 7124 5480
rect 6988 5104 7028 5144
rect 7180 5020 7220 5060
rect 6892 4936 6932 4976
rect 6796 4852 6836 4892
rect 6220 3676 6260 3716
rect 7276 4852 7316 4892
rect 7276 4096 7316 4136
rect 5644 3592 5684 3632
rect 6316 3592 6356 3632
rect 5452 3340 5492 3380
rect 5356 3088 5396 3128
rect 7660 6364 7700 6404
rect 7660 5440 7700 5480
rect 6316 3424 6356 3464
rect 5836 3256 5876 3296
rect 5356 2752 5396 2792
rect 3820 2500 3860 2540
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 3820 1912 3860 1952
rect 4396 1912 4436 1952
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 2956 1240 2996 1280
rect 4108 1240 4148 1280
rect 6508 3424 6548 3464
rect 6412 3256 6452 3296
rect 7084 3508 7124 3548
rect 7276 3508 7316 3548
rect 6988 3424 7028 3464
rect 7180 3340 7220 3380
rect 6700 3256 6740 3296
rect 6988 3256 7028 3296
rect 6604 2584 6644 2624
rect 6220 2500 6260 2540
rect 6796 2500 6836 2540
rect 7180 2500 7220 2540
rect 7468 3928 7508 3968
rect 8236 7960 8276 8000
rect 8716 7960 8756 8000
rect 8140 7876 8180 7916
rect 8044 7708 8084 7748
rect 9196 7876 9236 7916
rect 11404 10984 11444 11024
rect 12268 12328 12308 12368
rect 12076 12244 12116 12284
rect 11692 11656 11732 11696
rect 11692 11320 11732 11360
rect 11308 10732 11348 10772
rect 11020 10144 11060 10184
rect 10924 9388 10964 9428
rect 11212 9556 11252 9596
rect 11404 10144 11444 10184
rect 11788 10984 11828 11024
rect 12940 12328 12980 12368
rect 12364 12244 12404 12284
rect 12748 12244 12788 12284
rect 13132 11656 13172 11696
rect 11884 10732 11924 10772
rect 11500 9472 11540 9512
rect 11404 9388 11444 9428
rect 12172 9976 12212 10016
rect 11596 9388 11636 9428
rect 11884 9472 11924 9512
rect 12076 9472 12116 9512
rect 11884 9304 11924 9344
rect 11500 8800 11540 8840
rect 10156 7876 10196 7916
rect 9580 7288 9620 7328
rect 8524 7120 8564 7160
rect 8908 7120 8948 7160
rect 8812 7036 8852 7076
rect 9100 6364 9140 6404
rect 8140 5944 8180 5984
rect 8044 5608 8084 5648
rect 8812 5608 8852 5648
rect 8236 5440 8276 5480
rect 8716 4936 8756 4976
rect 9388 5860 9428 5900
rect 9196 5608 9236 5648
rect 7852 4096 7892 4136
rect 9100 4768 9140 4808
rect 9676 4768 9716 4808
rect 8908 4096 8948 4136
rect 7948 3928 7988 3968
rect 7756 3844 7796 3884
rect 7660 3508 7700 3548
rect 7948 3424 7988 3464
rect 7564 2584 7604 2624
rect 9388 3508 9428 3548
rect 8812 3424 8852 3464
rect 9388 3340 9428 3380
rect 8812 3256 8852 3296
rect 8620 3172 8660 3212
rect 9100 3172 9140 3212
rect 10636 7960 10676 8000
rect 10828 7960 10868 8000
rect 11308 7960 11348 8000
rect 12172 8800 12212 8840
rect 12748 9976 12788 10016
rect 12652 9472 12692 9512
rect 14284 11152 14324 11192
rect 13516 9556 13556 9596
rect 13804 9472 13844 9512
rect 13324 9304 13364 9344
rect 13708 9304 13748 9344
rect 12460 8044 12500 8084
rect 13516 7960 13556 8000
rect 10444 7540 10484 7580
rect 10444 6364 10484 6404
rect 11692 7540 11732 7580
rect 10924 7288 10964 7328
rect 10732 7120 10772 7160
rect 11788 7288 11828 7328
rect 11404 5944 11444 5984
rect 10828 4768 10868 4808
rect 7084 1912 7124 1952
rect 10348 4096 10388 4136
rect 10828 4012 10868 4052
rect 10732 3760 10772 3800
rect 10636 3424 10676 3464
rect 10924 3424 10964 3464
rect 10252 3256 10292 3296
rect 10060 2836 10100 2876
rect 10828 2836 10868 2876
rect 11788 4936 11828 4976
rect 11980 4852 12020 4892
rect 11212 4096 11252 4136
rect 11692 3928 11732 3968
rect 11212 3592 11252 3632
rect 11308 3508 11348 3548
rect 12076 4096 12116 4136
rect 12076 3928 12116 3968
rect 11884 3424 11924 3464
rect 13132 4936 13172 4976
rect 14284 8044 14324 8084
rect 12172 3592 12212 3632
rect 13132 3928 13172 3968
rect 13804 3760 13844 3800
rect 14284 3760 14324 3800
rect 12268 3424 12308 3464
rect 9964 2080 10004 2120
rect 10924 2080 10964 2120
rect 7084 1240 7124 1280
rect 7948 1240 7988 1280
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
<< metal3 >>
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 7363 13168 7372 13208
rect 7412 13168 8812 13208
rect 8852 13168 9484 13208
rect 9524 13168 9533 13208
rect 9091 13084 9100 13124
rect 9140 13084 10348 13124
rect 10388 13084 10924 13124
rect 10964 13084 10973 13124
rect 10531 13000 10540 13040
rect 10580 13000 11020 13040
rect 11060 13000 11692 13040
rect 11732 13000 11741 13040
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 7075 12832 7084 12872
rect 7124 12832 7852 12872
rect 7892 12832 8428 12872
rect 8468 12832 8908 12872
rect 8948 12832 8957 12872
rect 7363 12580 7372 12620
rect 7412 12580 9964 12620
rect 10004 12580 10013 12620
rect 10435 12580 10444 12620
rect 10484 12580 11500 12620
rect 11540 12580 11549 12620
rect 4099 12496 4108 12536
rect 4148 12496 4972 12536
rect 5012 12496 5021 12536
rect 7267 12496 7276 12536
rect 7316 12496 7564 12536
rect 7604 12496 7613 12536
rect 7171 12412 7180 12452
rect 7220 12412 7948 12452
rect 7988 12412 8812 12452
rect 8852 12412 8861 12452
rect 12259 12328 12268 12368
rect 12308 12328 12940 12368
rect 12980 12328 12989 12368
rect 2179 12244 2188 12284
rect 2228 12244 2764 12284
rect 2804 12244 2813 12284
rect 4771 12244 4780 12284
rect 4820 12244 5260 12284
rect 5300 12244 5309 12284
rect 12067 12244 12076 12284
rect 12116 12244 12364 12284
rect 12404 12244 12748 12284
rect 12788 12244 12797 12284
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 8707 11824 8716 11864
rect 8756 11824 9100 11864
rect 9140 11824 10060 11864
rect 10100 11824 10109 11864
rect 3331 11656 3340 11696
rect 3380 11656 4108 11696
rect 4148 11656 4157 11696
rect 6307 11656 6316 11696
rect 6356 11656 7276 11696
rect 7316 11656 7325 11696
rect 9955 11656 9964 11696
rect 10004 11656 11692 11696
rect 11732 11656 13132 11696
rect 13172 11656 13181 11696
rect 7459 11404 7468 11444
rect 7508 11404 8908 11444
rect 8948 11404 8957 11444
rect 9859 11404 9868 11444
rect 9908 11404 10156 11444
rect 10196 11404 10205 11444
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 7555 11320 7564 11360
rect 7604 11320 8716 11360
rect 8756 11320 9964 11360
rect 10004 11320 10013 11360
rect 10435 11320 10444 11360
rect 10484 11320 11692 11360
rect 11732 11320 11741 11360
rect 0 11192 80 11212
rect 14920 11192 15000 11212
rect 0 11152 844 11192
rect 884 11152 893 11192
rect 14275 11152 14284 11192
rect 14324 11152 15000 11192
rect 0 11132 80 11152
rect 14920 11132 15000 11152
rect 7459 11068 7468 11108
rect 7508 11068 9004 11108
rect 9044 11068 9053 11108
rect 1891 10984 1900 11024
rect 1940 10984 3436 11024
rect 3476 10984 4204 11024
rect 4244 10984 4492 11024
rect 4532 10984 4541 11024
rect 6883 10984 6892 11024
rect 6932 10984 7852 11024
rect 7892 10984 7901 11024
rect 11395 10984 11404 11024
rect 11444 10984 11788 11024
rect 11828 10984 11837 11024
rect 9571 10732 9580 10772
rect 9620 10732 10540 10772
rect 10580 10732 10732 10772
rect 10772 10732 11308 10772
rect 11348 10732 11884 10772
rect 11924 10732 11933 10772
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 4483 10396 4492 10436
rect 4532 10396 5260 10436
rect 5300 10396 5309 10436
rect 6115 10312 6124 10352
rect 6164 10312 7276 10352
rect 7316 10312 7325 10352
rect 9859 10312 9868 10352
rect 9908 10312 10292 10352
rect 10252 10268 10292 10312
rect 9580 10228 10060 10268
rect 10100 10228 10109 10268
rect 10243 10228 10252 10268
rect 10292 10228 10636 10268
rect 10676 10228 10685 10268
rect 6019 10144 6028 10184
rect 6068 10144 6892 10184
rect 6932 10144 6941 10184
rect 8995 10144 9004 10184
rect 9044 10144 9484 10184
rect 9524 10144 9533 10184
rect 9580 10100 9620 10228
rect 9763 10144 9772 10184
rect 9812 10144 10348 10184
rect 10388 10144 10732 10184
rect 10772 10144 10781 10184
rect 11011 10144 11020 10184
rect 11060 10144 11404 10184
rect 11444 10144 11453 10184
rect 8131 10060 8140 10100
rect 8180 10060 9620 10100
rect 9667 10060 9676 10100
rect 9716 10060 10156 10100
rect 10196 10060 10205 10100
rect 9475 9976 9484 10016
rect 9524 9976 10060 10016
rect 10100 9976 10109 10016
rect 12163 9976 12172 10016
rect 12212 9976 12748 10016
rect 12788 9976 12797 10016
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 11203 9556 11212 9596
rect 11252 9556 13516 9596
rect 13556 9556 13565 9596
rect 11491 9472 11500 9512
rect 11540 9472 11884 9512
rect 11924 9472 11933 9512
rect 12067 9472 12076 9512
rect 12116 9472 12652 9512
rect 12692 9472 12701 9512
rect 13795 9472 13804 9512
rect 13844 9472 13853 9512
rect 13804 9428 13844 9472
rect 10339 9388 10348 9428
rect 10388 9388 10924 9428
rect 10964 9388 10973 9428
rect 11395 9388 11404 9428
rect 11444 9388 11596 9428
rect 11636 9388 13844 9428
rect 11875 9304 11884 9344
rect 11924 9304 13324 9344
rect 13364 9304 13708 9344
rect 13748 9304 13757 9344
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 8515 8800 8524 8840
rect 8564 8800 9388 8840
rect 9428 8800 9437 8840
rect 11491 8800 11500 8840
rect 11540 8800 12172 8840
rect 12212 8800 12221 8840
rect 3331 8632 3340 8672
rect 3380 8632 3724 8672
rect 3764 8632 3773 8672
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 12451 8044 12460 8084
rect 12500 8044 14284 8084
rect 14324 8044 14333 8084
rect 3235 7960 3244 8000
rect 3284 7960 4396 8000
rect 4436 7960 4445 8000
rect 4675 7960 4684 8000
rect 4724 7960 5740 8000
rect 5780 7960 5789 8000
rect 7459 7960 7468 8000
rect 7508 7960 8236 8000
rect 8276 7960 8285 8000
rect 8707 7960 8716 8000
rect 8756 7960 10636 8000
rect 10676 7960 10828 8000
rect 10868 7960 10877 8000
rect 11299 7960 11308 8000
rect 11348 7960 13516 8000
rect 13556 7960 13565 8000
rect 8131 7876 8140 7916
rect 8180 7876 9196 7916
rect 9236 7876 10156 7916
rect 10196 7876 10205 7916
rect 3331 7792 3340 7832
rect 3380 7792 4204 7832
rect 4244 7792 4253 7832
rect 5539 7792 5548 7832
rect 5588 7792 6796 7832
rect 6836 7792 6845 7832
rect 1123 7708 1132 7748
rect 1172 7708 2188 7748
rect 2228 7708 2237 7748
rect 4867 7708 4876 7748
rect 4916 7708 8044 7748
rect 8084 7708 8093 7748
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 10435 7540 10444 7580
rect 10484 7540 11692 7580
rect 11732 7540 11741 7580
rect 4771 7372 4780 7412
rect 4820 7372 4972 7412
rect 5012 7372 5021 7412
rect 9571 7288 9580 7328
rect 9620 7288 9629 7328
rect 10915 7288 10924 7328
rect 10964 7288 11788 7328
rect 11828 7288 11837 7328
rect 6019 7204 6028 7244
rect 6068 7204 6604 7244
rect 6644 7204 6653 7244
rect 9580 7160 9620 7288
rect 4771 7120 4780 7160
rect 4820 7120 5452 7160
rect 5492 7120 5501 7160
rect 5923 7120 5932 7160
rect 5972 7120 6508 7160
rect 6548 7120 6557 7160
rect 7555 7120 7564 7160
rect 7604 7120 8524 7160
rect 8564 7120 8573 7160
rect 8899 7120 8908 7160
rect 8948 7120 10732 7160
rect 10772 7120 10781 7160
rect 7459 7036 7468 7076
rect 7508 7036 8812 7076
rect 8852 7036 8861 7076
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 3523 6700 3532 6740
rect 3572 6700 4012 6740
rect 4052 6700 6320 6740
rect 6280 6572 6320 6700
rect 6280 6532 6508 6572
rect 6548 6532 6557 6572
rect 2659 6448 2668 6488
rect 2708 6448 4108 6488
rect 4148 6448 4157 6488
rect 5539 6448 5548 6488
rect 5588 6448 6028 6488
rect 6068 6448 6077 6488
rect 6211 6448 6220 6488
rect 6260 6448 7276 6488
rect 7316 6448 7325 6488
rect 5155 6364 5164 6404
rect 5204 6364 7372 6404
rect 7412 6364 7421 6404
rect 7651 6364 7660 6404
rect 7700 6364 9100 6404
rect 9140 6364 10444 6404
rect 10484 6364 10493 6404
rect 5028 6280 5068 6320
rect 5108 6280 5117 6320
rect 5700 6280 5740 6320
rect 5780 6280 5789 6320
rect 6028 6280 6316 6320
rect 6356 6280 6365 6320
rect 5068 6236 5108 6280
rect 5740 6236 5780 6280
rect 6028 6236 6068 6280
rect 5068 6196 6068 6236
rect 6115 6196 6124 6236
rect 6164 6196 6796 6236
rect 6836 6196 6845 6236
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 8131 5944 8140 5984
rect 8180 5944 11404 5984
rect 11444 5944 11453 5984
rect 7267 5860 7276 5900
rect 7316 5860 9388 5900
rect 9428 5860 9437 5900
rect 4771 5692 4780 5732
rect 4820 5692 4972 5732
rect 5012 5692 5644 5732
rect 5684 5692 6508 5732
rect 6548 5692 6557 5732
rect 4675 5608 4684 5648
rect 4724 5608 5068 5648
rect 5108 5608 5932 5648
rect 5972 5608 5981 5648
rect 6595 5608 6604 5648
rect 6644 5608 8044 5648
rect 8084 5608 8093 5648
rect 8803 5608 8812 5648
rect 8852 5608 9196 5648
rect 9236 5608 9245 5648
rect 4483 5440 4492 5480
rect 4532 5440 5836 5480
rect 5876 5440 6220 5480
rect 6260 5440 6269 5480
rect 6499 5440 6508 5480
rect 6548 5440 7084 5480
rect 7124 5440 7133 5480
rect 7651 5440 7660 5480
rect 7700 5440 8236 5480
rect 8276 5440 8285 5480
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 5155 5104 5164 5144
rect 5204 5104 6988 5144
rect 7028 5104 7037 5144
rect 1987 5020 1996 5060
rect 2036 5020 3724 5060
rect 3764 5020 3773 5060
rect 6691 5020 6700 5060
rect 6740 5020 7180 5060
rect 7220 5020 7229 5060
rect 2179 4936 2188 4976
rect 2228 4936 2380 4976
rect 2420 4936 4012 4976
rect 4052 4936 4061 4976
rect 4291 4936 4300 4976
rect 4340 4936 5452 4976
rect 5492 4936 5501 4976
rect 6499 4936 6508 4976
rect 6548 4936 6892 4976
rect 6932 4936 8716 4976
rect 8756 4936 8765 4976
rect 11779 4936 11788 4976
rect 11828 4936 13132 4976
rect 13172 4936 13181 4976
rect 6787 4852 6796 4892
rect 6836 4852 7276 4892
rect 7316 4852 11980 4892
rect 12020 4852 12029 4892
rect 9091 4768 9100 4808
rect 9140 4768 9676 4808
rect 9716 4768 10828 4808
rect 10868 4768 10877 4808
rect 3907 4684 3916 4724
rect 3956 4684 4492 4724
rect 4532 4684 4972 4724
rect 5012 4684 5356 4724
rect 5396 4684 5405 4724
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 931 4348 940 4388
rect 980 4348 1612 4388
rect 1652 4348 1661 4388
rect 1699 4096 1708 4136
rect 1748 4096 2668 4136
rect 2708 4096 4300 4136
rect 4340 4096 5548 4136
rect 5588 4096 5597 4136
rect 7267 4096 7276 4136
rect 7316 4096 7852 4136
rect 7892 4096 8908 4136
rect 8948 4096 8957 4136
rect 10339 4096 10348 4136
rect 10388 4096 11212 4136
rect 11252 4096 11261 4136
rect 12067 4096 12076 4136
rect 12116 4096 12125 4136
rect 12076 4052 12116 4096
rect 10819 4012 10828 4052
rect 10868 4012 12116 4052
rect 7459 3928 7468 3968
rect 7508 3928 7948 3968
rect 7988 3928 7997 3968
rect 11683 3928 11692 3968
rect 11732 3928 12076 3968
rect 12116 3928 13132 3968
rect 13172 3928 13181 3968
rect 2284 3844 7756 3884
rect 7796 3844 7805 3884
rect 0 3800 80 3820
rect 2284 3800 2324 3844
rect 14920 3800 15000 3820
rect 0 3760 2324 3800
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 4867 3760 4876 3800
rect 4916 3760 5164 3800
rect 5204 3760 5213 3800
rect 10723 3760 10732 3800
rect 10772 3760 13804 3800
rect 13844 3760 13853 3800
rect 14275 3760 14284 3800
rect 14324 3760 15000 3800
rect 0 3740 80 3760
rect 14920 3740 15000 3760
rect 4771 3676 4780 3716
rect 4820 3676 6220 3716
rect 6260 3676 6269 3716
rect 5059 3592 5068 3632
rect 5108 3592 5644 3632
rect 5684 3592 5693 3632
rect 6280 3592 6316 3632
rect 6356 3592 6365 3632
rect 11203 3592 11212 3632
rect 11252 3592 12172 3632
rect 12212 3592 12221 3632
rect 6280 3548 6320 3592
rect 2659 3508 2668 3548
rect 2708 3508 6320 3548
rect 7075 3508 7084 3548
rect 7124 3508 7276 3548
rect 7316 3508 7660 3548
rect 7700 3508 9388 3548
rect 9428 3508 9437 3548
rect 10636 3508 11308 3548
rect 11348 3508 11357 3548
rect 10636 3464 10676 3508
rect 2467 3424 2476 3464
rect 2516 3424 3052 3464
rect 3092 3424 3101 3464
rect 6307 3424 6316 3464
rect 6356 3424 6508 3464
rect 6548 3424 6557 3464
rect 6979 3424 6988 3464
rect 7028 3424 7948 3464
rect 7988 3424 7997 3464
rect 8803 3424 8812 3464
rect 8852 3424 10636 3464
rect 10676 3424 10685 3464
rect 10915 3424 10924 3464
rect 10964 3424 11884 3464
rect 11924 3424 12268 3464
rect 12308 3424 12317 3464
rect 4387 3340 4396 3380
rect 4436 3340 4876 3380
rect 4916 3340 5452 3380
rect 5492 3340 5501 3380
rect 7171 3340 7180 3380
rect 7220 3340 9388 3380
rect 9428 3340 9437 3380
rect 5827 3256 5836 3296
rect 5876 3256 6412 3296
rect 6452 3256 6700 3296
rect 6740 3256 6988 3296
rect 7028 3256 7037 3296
rect 8803 3256 8812 3296
rect 8852 3256 10252 3296
rect 10292 3256 10301 3296
rect 8611 3172 8620 3212
rect 8660 3172 9100 3212
rect 9140 3172 9149 3212
rect 4867 3088 4876 3128
rect 4916 3088 5356 3128
rect 5396 3088 5405 3128
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 10051 2836 10060 2876
rect 10100 2836 10828 2876
rect 10868 2836 10877 2876
rect 4771 2752 4780 2792
rect 4820 2752 5356 2792
rect 5396 2752 5405 2792
rect 6595 2584 6604 2624
rect 6644 2584 7564 2624
rect 7604 2584 7613 2624
rect 3235 2500 3244 2540
rect 3284 2500 3820 2540
rect 3860 2500 3869 2540
rect 6211 2500 6220 2540
rect 6260 2500 6796 2540
rect 6836 2500 7180 2540
rect 7220 2500 7229 2540
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 9955 2080 9964 2120
rect 10004 2080 10924 2120
rect 10964 2080 10973 2120
rect 3811 1912 3820 1952
rect 3860 1912 4396 1952
rect 4436 1912 7084 1952
rect 7124 1912 7133 1952
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 2947 1240 2956 1280
rect 2996 1240 4108 1280
rect 4148 1240 4157 1280
rect 7075 1240 7084 1280
rect 7124 1240 7948 1280
rect 7988 1240 7997 1280
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
<< via3 >>
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
<< metal4 >>
rect 3076 13628 3516 13652
rect 3076 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3516 13628
rect 3076 12116 3516 13588
rect 3076 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3516 12116
rect 3076 10604 3516 12076
rect 3076 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3516 10604
rect 3076 9092 3516 10564
rect 3076 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3516 9092
rect 3076 7580 3516 9052
rect 3076 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3516 7580
rect 3076 6068 3516 7540
rect 3076 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3516 6068
rect 3076 4556 3516 6028
rect 3076 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3516 4556
rect 3076 3640 3516 4516
rect 3076 3600 3132 3640
rect 3172 3600 3228 3640
rect 3268 3600 3324 3640
rect 3364 3600 3420 3640
rect 3460 3600 3516 3640
rect 3076 3544 3516 3600
rect 3076 3504 3132 3544
rect 3172 3504 3228 3544
rect 3268 3504 3324 3544
rect 3364 3504 3420 3544
rect 3460 3504 3516 3544
rect 3076 3448 3516 3504
rect 3076 3408 3132 3448
rect 3172 3408 3228 3448
rect 3268 3408 3324 3448
rect 3364 3408 3420 3448
rect 3460 3408 3516 3448
rect 3076 3352 3516 3408
rect 3076 3312 3132 3352
rect 3172 3312 3228 3352
rect 3268 3312 3324 3352
rect 3364 3312 3420 3352
rect 3460 3312 3516 3352
rect 3076 3044 3516 3312
rect 3076 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3516 3044
rect 3076 1532 3516 3004
rect 3076 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3516 1532
rect 3076 712 3516 1492
rect 4316 12872 4756 13652
rect 4316 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4756 12872
rect 4316 11360 4756 12832
rect 4316 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4756 11360
rect 4316 9848 4756 11320
rect 4316 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4756 9848
rect 4316 8336 4756 9808
rect 4316 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4756 8336
rect 4316 6824 4756 8296
rect 4316 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4756 6824
rect 4316 5312 4756 6784
rect 4316 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4756 5312
rect 4316 4880 4756 5272
rect 4316 4840 4372 4880
rect 4412 4840 4468 4880
rect 4508 4840 4564 4880
rect 4604 4840 4660 4880
rect 4700 4840 4756 4880
rect 4316 4784 4756 4840
rect 4316 4744 4372 4784
rect 4412 4744 4468 4784
rect 4508 4744 4564 4784
rect 4604 4744 4660 4784
rect 4700 4744 4756 4784
rect 4316 4688 4756 4744
rect 4316 4648 4372 4688
rect 4412 4648 4468 4688
rect 4508 4648 4564 4688
rect 4604 4648 4660 4688
rect 4700 4648 4756 4688
rect 4316 4592 4756 4648
rect 4316 4552 4372 4592
rect 4412 4552 4468 4592
rect 4508 4552 4564 4592
rect 4604 4552 4660 4592
rect 4700 4552 4756 4592
rect 4316 3800 4756 4552
rect 4316 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4756 3800
rect 4316 2288 4756 3760
rect 4316 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4756 2288
rect 4316 776 4756 2248
rect 4316 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4756 776
rect 4316 712 4756 736
<< via4 >>
rect 3132 3600 3172 3640
rect 3228 3600 3268 3640
rect 3324 3600 3364 3640
rect 3420 3600 3460 3640
rect 3132 3504 3172 3544
rect 3228 3504 3268 3544
rect 3324 3504 3364 3544
rect 3420 3504 3460 3544
rect 3132 3408 3172 3448
rect 3228 3408 3268 3448
rect 3324 3408 3364 3448
rect 3420 3408 3460 3448
rect 3132 3312 3172 3352
rect 3228 3312 3268 3352
rect 3324 3312 3364 3352
rect 3420 3312 3460 3352
rect 4372 4840 4412 4880
rect 4468 4840 4508 4880
rect 4564 4840 4604 4880
rect 4660 4840 4700 4880
rect 4372 4744 4412 4784
rect 4468 4744 4508 4784
rect 4564 4744 4604 4784
rect 4660 4744 4700 4784
rect 4372 4648 4412 4688
rect 4468 4648 4508 4688
rect 4564 4648 4604 4688
rect 4660 4648 4700 4688
rect 4372 4552 4412 4592
rect 4468 4552 4508 4592
rect 4564 4552 4604 4592
rect 4660 4552 4700 4592
<< metal5 >>
rect 532 4880 14444 4936
rect 532 4840 4372 4880
rect 4412 4840 4468 4880
rect 4508 4840 4564 4880
rect 4604 4840 4660 4880
rect 4700 4840 14444 4880
rect 532 4784 14444 4840
rect 532 4744 4372 4784
rect 4412 4744 4468 4784
rect 4508 4744 4564 4784
rect 4604 4744 4660 4784
rect 4700 4744 14444 4784
rect 532 4688 14444 4744
rect 532 4648 4372 4688
rect 4412 4648 4468 4688
rect 4508 4648 4564 4688
rect 4604 4648 4660 4688
rect 4700 4648 14444 4688
rect 532 4592 14444 4648
rect 532 4552 4372 4592
rect 4412 4552 4468 4592
rect 4508 4552 4564 4592
rect 4604 4552 4660 4592
rect 4700 4552 14444 4592
rect 532 4496 14444 4552
rect 532 3640 14444 3696
rect 532 3600 3132 3640
rect 3172 3600 3228 3640
rect 3268 3600 3324 3640
rect 3364 3600 3420 3640
rect 3460 3600 14444 3640
rect 532 3544 14444 3600
rect 532 3504 3132 3544
rect 3172 3504 3228 3544
rect 3268 3504 3324 3544
rect 3364 3504 3420 3544
rect 3460 3504 14444 3544
rect 532 3448 14444 3504
rect 532 3408 3132 3448
rect 3172 3408 3228 3448
rect 3268 3408 3324 3448
rect 3364 3408 3420 3448
rect 3460 3408 14444 3448
rect 532 3352 14444 3408
rect 532 3312 3132 3352
rect 3172 3312 3228 3352
rect 3268 3312 3324 3352
rect 3364 3312 3420 3352
rect 3460 3312 14444 3352
rect 532 3256 14444 3312
use sg13g2_inv_1  _082_
timestamp 1676382929
transform -1 0 1824 0 1 3780
box -48 -56 336 834
use sg13g2_inv_1  _083_
timestamp 1676382929
transform -1 0 6336 0 -1 6804
box -48 -56 336 834
use sg13g2_inv_1  _084_
timestamp 1676382929
transform -1 0 5760 0 1 8316
box -48 -56 336 834
use sg13g2_nand3_1  _085_
timestamp 1683988354
transform -1 0 5184 0 1 2268
box -48 -56 528 834
use sg13g2_and4_1  _086_
timestamp 1676985977
transform 1 0 5184 0 -1 3780
box -48 -56 816 834
use sg13g2_and2_1  _087_
timestamp 1676901763
transform 1 0 6336 0 1 3780
box -48 -56 528 834
use sg13g2_nand4_1  _088_
timestamp 1685201930
transform 1 0 6912 0 1 2268
box -48 -56 624 834
use sg13g2_nor2_1  _089_
timestamp 1676627187
transform 1 0 8640 0 1 3780
box -48 -56 432 834
use sg13g2_nand2_1  _090_
timestamp 1676557249
transform -1 0 12192 0 -1 3780
box -48 -56 432 834
use sg13g2_nor3_1  _091_
timestamp 1676639442
transform 1 0 6432 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _092_
timestamp 1676557249
transform -1 0 9024 0 1 6804
box -48 -56 432 834
use sg13g2_nor4_2  _093_
timestamp 1685199459
transform 1 0 6624 0 1 5292
box -48 -56 1200 834
use sg13g2_nand3_1  _094_
timestamp 1683988354
transform -1 0 4896 0 1 5292
box -48 -56 528 834
use sg13g2_nand4_1  _095_
timestamp 1685201930
transform -1 0 6624 0 1 5292
box -48 -56 624 834
use sg13g2_nor2_1  _096_
timestamp 1676627187
transform 1 0 5184 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2b_1  _097_
timestamp 1685181386
transform 1 0 4896 0 -1 12852
box -54 -56 528 834
use sg13g2_xor2_1  _098_
timestamp 1677577977
transform 1 0 11712 0 -1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _099_
timestamp 1677516600
transform 1 0 9792 0 1 11340
box -48 -56 816 834
use sg13g2_xnor2_1  _100_
timestamp 1677516600
transform -1 0 12288 0 1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _101_
timestamp 1685175443
transform -1 0 11616 0 -1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _102_
timestamp 1683973020
transform 1 0 13440 0 -1 9828
box -48 -56 528 834
use sg13g2_xor2_1  _103_
timestamp 1677577977
transform -1 0 11712 0 -1 8316
box -48 -56 816 834
use sg13g2_xnor2_1  _104_
timestamp 1677516600
transform -1 0 8352 0 -1 12852
box -48 -56 816 834
use sg13g2_nor2_1  _105_
timestamp 1676627187
transform -1 0 7584 0 -1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _106_
timestamp 1683973020
transform -1 0 7488 0 1 12852
box -48 -56 528 834
use sg13g2_and3_1  _107_
timestamp 1676971669
transform 1 0 8544 0 1 12852
box -48 -56 720 834
use sg13g2_nor3_1  _108_
timestamp 1676639442
transform 1 0 8928 0 1 9828
box -48 -56 528 834
use sg13g2_nor2_1  _109_
timestamp 1676627187
transform -1 0 10656 0 1 12852
box -48 -56 432 834
use sg13g2_and2_1  _110_
timestamp 1676901763
transform -1 0 11136 0 1 12852
box -48 -56 528 834
use sg13g2_nor3_1  _111_
timestamp 1676639442
transform -1 0 10656 0 1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  _112_
timestamp 1683973020
transform 1 0 9504 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _113_
timestamp 1685175443
transform -1 0 10464 0 1 9828
box -48 -56 538 834
use sg13g2_inv_1  _114_
timestamp 1676382929
transform -1 0 9600 0 1 8316
box -48 -56 336 834
use sg13g2_xor2_1  _115_
timestamp 1677577977
transform -1 0 4416 0 -1 5292
box -48 -56 816 834
use sg13g2_a21o_1  _116_
timestamp 1677175127
transform -1 0 5952 0 -1 5292
box -48 -56 720 834
use sg13g2_and2_1  _117_
timestamp 1676901763
transform 1 0 5952 0 -1 5292
box -48 -56 528 834
use sg13g2_xnor2_1  _118_
timestamp 1677516600
transform -1 0 5664 0 1 756
box -48 -56 816 834
use sg13g2_xor2_1  _119_
timestamp 1677577977
transform 1 0 6048 0 -1 3780
box -48 -56 816 834
use sg13g2_xor2_1  _120_
timestamp 1677577977
transform 1 0 7584 0 -1 3780
box -48 -56 816 834
use sg13g2_a21o_1  _121_
timestamp 1677175127
transform -1 0 7584 0 -1 3780
box -48 -56 720 834
use sg13g2_and2_1  _122_
timestamp 1676901763
transform 1 0 7776 0 1 3780
box -48 -56 528 834
use sg13g2_xnor2_1  _123_
timestamp 1677516600
transform 1 0 7008 0 1 3780
box -48 -56 816 834
use sg13g2_xor2_1  _124_
timestamp 1677577977
transform -1 0 11808 0 -1 3780
box -48 -56 816 834
use sg13g2_a21oi_1  _125_
timestamp 1683973020
transform -1 0 11040 0 -1 3780
box -48 -56 528 834
use sg13g2_nor2_1  _126_
timestamp 1676627187
transform 1 0 10080 0 -1 8316
box -48 -56 432 834
use sg13g2_xor2_1  _127_
timestamp 1677577977
transform -1 0 9696 0 -1 8316
box -48 -56 816 834
use sg13g2_a21oi_1  _128_
timestamp 1683973020
transform -1 0 8448 0 1 5292
box -48 -56 528 834
use sg13g2_nor2_1  _129_
timestamp 1676627187
transform 1 0 4896 0 1 5292
box -48 -56 432 834
use sg13g2_xor2_1  _130_
timestamp 1677577977
transform -1 0 6048 0 1 5292
box -48 -56 816 834
use sg13g2_a21o_1  _131_
timestamp 1677175127
transform 1 0 4320 0 -1 8316
box -48 -56 720 834
use sg13g2_and2_1  _132_
timestamp 1676901763
transform -1 0 3456 0 -1 8316
box -48 -56 528 834
use sg13g2_xnor2_1  _133_
timestamp 1677516600
transform -1 0 3648 0 -1 9828
box -48 -56 816 834
use sg13g2_xnor2_1  _134_
timestamp 1677516600
transform 1 0 5280 0 -1 6804
box -48 -56 816 834
use sg13g2_mux2_1  _135_
timestamp 1677247768
transform 1 0 11616 0 -1 9828
box -48 -56 1008 834
use sg13g2_tiehi  _136__6
timestamp 1680000651
transform -1 0 12672 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_2  _136_
timestamp 1746535184
transform 1 0 11712 0 1 8316
box -48 -56 2736 834
use sg13g2_tiehi  _137__7
timestamp 1680000651
transform -1 0 1440 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _137_
timestamp 1746535128
transform 1 0 576 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _138__8
timestamp 1680000651
transform 1 0 2304 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _138_
timestamp 1746535128
transform 1 0 2112 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _139__9
timestamp 1680000651
transform -1 0 4032 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _139_
timestamp 1746535128
transform 1 0 3264 0 1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _140__31
timestamp 1680000651
transform -1 0 5568 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _140_
timestamp 1746535128
transform 1 0 4704 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _141__5
timestamp 1680000651
transform -1 0 7584 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_2  _141_
timestamp 1746535184
transform 1 0 5568 0 -1 9828
box -48 -56 2736 834
use sg13g2_tiehi  _142__20
timestamp 1680000651
transform -1 0 7104 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_2  _142_
timestamp 1746535184
transform 1 0 6240 0 1 11340
box -48 -56 2736 834
use sg13g2_tiehi  _143__18
timestamp 1680000651
transform 1 0 6624 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _143_
timestamp 1746535128
transform 1 0 7392 0 -1 11340
box -48 -56 2640 834
use sg13g2_tiehi  _144__16
timestamp 1680000651
transform -1 0 11520 0 1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _144_
timestamp 1746535128
transform 1 0 10272 0 -1 12852
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _145_
timestamp 1746535128
transform 1 0 8448 0 -1 9828
box -48 -56 2640 834
use sg13g2_tiehi  _145__14
timestamp 1680000651
transform -1 0 9312 0 1 8316
box -48 -56 432 834
use sg13g2_tiehi  _146__12
timestamp 1680000651
transform -1 0 1728 0 1 5292
box -48 -56 432 834
use sg13g2_dfrbpq_2  _146_
timestamp 1746535184
transform 1 0 864 0 -1 5292
box -48 -56 2736 834
use sg13g2_tiehi  _147__11
timestamp 1680000651
transform 1 0 1824 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _147_
timestamp 1746535128
transform 1 0 1920 0 1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _148__10
timestamp 1680000651
transform 1 0 2208 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _148_
timestamp 1746535128
transform 1 0 2592 0 -1 3780
box -48 -56 2640 834
use sg13g2_tiehi  _149__4
timestamp 1680000651
transform -1 0 3936 0 1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _149_
timestamp 1746535128
transform 1 0 3072 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _150__30
timestamp 1680000651
transform 1 0 6816 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _150_
timestamp 1746535128
transform -1 0 8448 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _151__29
timestamp 1680000651
transform -1 0 9696 0 1 756
box -48 -56 432 834
use sg13g2_dfrbpq_1  _151_
timestamp 1746535128
transform 1 0 8448 0 -1 2268
box -48 -56 2640 834
use sg13g2_tiehi  _152__28
timestamp 1680000651
transform -1 0 10560 0 -1 3780
box -48 -56 432 834
use sg13g2_dfrbpq_1  _152_
timestamp 1746535128
transform 1 0 8352 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _153_
timestamp 1746535128
transform 1 0 7776 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _153__27
timestamp 1680000651
transform -1 0 8640 0 1 3780
box -48 -56 432 834
use sg13g2_tiehi  _154__26
timestamp 1680000651
transform -1 0 13056 0 -1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _154_
timestamp 1746535128
transform 1 0 11808 0 -1 5292
box -48 -56 2640 834
use sg13g2_tiehi  _155__25
timestamp 1680000651
transform -1 0 12096 0 1 6804
box -48 -56 432 834
use sg13g2_dfrbpq_1  _155_
timestamp 1746535128
transform 1 0 10464 0 1 5292
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _156_
timestamp 1746535128
transform 1 0 9120 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _156__24
timestamp 1680000651
transform -1 0 10368 0 -1 6804
box -48 -56 432 834
use sg13g2_tiehi  _157__23
timestamp 1680000651
transform -1 0 7200 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _157_
timestamp 1746535128
transform 1 0 6336 0 -1 6804
box -48 -56 2640 834
use sg13g2_dfrbpq_2  _158_
timestamp 1746535184
transform 1 0 2592 0 -1 6804
box -48 -56 2736 834
use sg13g2_tiehi  _158__22
timestamp 1680000651
transform -1 0 3456 0 1 5292
box -48 -56 432 834
use sg13g2_tiehi  _159__21
timestamp 1680000651
transform -1 0 4032 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _159_
timestamp 1746535128
transform 1 0 2880 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _160__19
timestamp 1680000651
transform -1 0 1920 0 -1 8316
box -48 -56 432 834
use sg13g2_dfrbpq_1  _160_
timestamp 1746535128
transform 1 0 1056 0 1 6804
box -48 -56 2640 834
use sg13g2_tiehi  _161__17
timestamp 1680000651
transform -1 0 6624 0 1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _161_
timestamp 1746535128
transform 1 0 5760 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _162__13
timestamp 1680000651
transform -1 0 14304 0 -1 9828
box -48 -56 432 834
use sg13g2_dfrbpq_1  _162_
timestamp 1746535128
transform -1 0 14400 0 -1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _163__15
timestamp 1680000651
transform -1 0 13248 0 -1 12852
box -48 -56 432 834
use sg13g2_dfrbpq_1  _163_
timestamp 1746535128
transform 1 0 11808 0 1 11340
box -48 -56 2640 834
use sg13g2_buf_8  clkbuf_0_clk
timestamp 1676451365
transform 1 0 7584 0 -1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_0__f_clk
timestamp 1676451365
transform -1 0 5184 0 1 3780
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_1__f_clk
timestamp 1676451365
transform 1 0 4800 0 1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_2__f_clk
timestamp 1676451365
transform 1 0 10368 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_2_3__f_clk
timestamp 1676451365
transform 1 0 10560 0 1 11340
box -48 -56 1296 834
use sg13g2_buf_1  clkload0
timestamp 1676381911
transform 1 0 4416 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  clkload1
timestamp 1676381911
transform 1 0 10944 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_35
timestamp 1677579658
transform 1 0 3936 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_53
timestamp 1679581782
transform 1 0 5664 0 1 756
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_60
timestamp 1679577901
transform 1 0 6336 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_64
timestamp 1677579658
transform 1 0 6720 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_69
timestamp 1679581782
transform 1 0 7200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_76
timestamp 1679581782
transform 1 0 7872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_83
timestamp 1679581782
transform 1 0 8544 0 1 756
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_90
timestamp 1677579658
transform 1 0 9216 0 1 756
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_95
timestamp 1679581782
transform 1 0 9696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_102
timestamp 1679581782
transform 1 0 10368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_109
timestamp 1679581782
transform 1 0 11040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_116
timestamp 1679581782
transform 1 0 11712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_123
timestamp 1679581782
transform 1 0 12384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_130
timestamp 1679581782
transform 1 0 13056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_137
timestamp 1679581782
transform 1 0 13728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_21
timestamp 1679577901
transform 1 0 2592 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_25
timestamp 1677579658
transform 1 0 2976 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_53
timestamp 1677580104
transform 1 0 5664 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_109
timestamp 1679581782
transform 1 0 11040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_116
timestamp 1679581782
transform 1 0 11712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_123
timestamp 1679581782
transform 1 0 12384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_130
timestamp 1679581782
transform 1 0 13056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_137
timestamp 1679581782
transform 1 0 13728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1248 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_41
timestamp 1677580104
transform 1 0 4512 0 1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 11328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 12000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 12672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679581782
transform 1 0 13344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_140
timestamp 1679577901
transform 1 0 14016 0 1 2268
box -48 -56 432 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 1920 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_56
timestamp 1677579658
transform 1 0 5952 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_65
timestamp 1677579658
transform 1 0 6816 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_90
timestamp 1677579658
transform 1 0 9216 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_121
timestamp 1679581782
transform 1 0 12192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_128
timestamp 1679581782
transform 1 0 12864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_135
timestamp 1679581782
transform 1 0 13536 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_142
timestamp 1677580104
transform 1 0 14208 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 576 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_7
timestamp 1677580104
transform 1 0 1248 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_9
timestamp 1677579658
transform 1 0 1440 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_30
timestamp 1677579658
transform 1 0 3456 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_48
timestamp 1677580104
transform 1 0 5184 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_59
timestamp 1677579658
transform 1 0 6240 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_65
timestamp 1677580104
transform 1 0 6816 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_88
timestamp 1677580104
transform 1 0 9024 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_90
timestamp 1677579658
transform 1 0 9216 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_100
timestamp 1677580104
transform 1 0 10176 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_102
timestamp 1677579658
transform 1 0 10368 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_139
timestamp 1677579658
transform 1 0 13920 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_0
timestamp 1677580104
transform 1 0 576 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_2
timestamp 1677579658
transform 1 0 768 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_31
timestamp 1677579658
transform 1 0 3552 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_115
timestamp 1677580104
transform 1 0 11616 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 576 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_7
timestamp 1677579658
transform 1 0 1248 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_12
timestamp 1679581782
transform 1 0 1728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_19
timestamp 1679581782
transform 1 0 2400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_30
timestamp 1679581782
transform 1 0 3456 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_37
timestamp 1677580104
transform 1 0 4128 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_39
timestamp 1677579658
transform 1 0 4320 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_75
timestamp 1677580104
transform 1 0 7776 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_100
timestamp 1677580104
transform 1 0 10176 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_102
timestamp 1677579658
transform 1 0 10368 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_130
timestamp 1679581782
transform 1 0 13056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_137
timestamp 1679581782
transform 1 0 13728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 1920 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_87
timestamp 1677580104
transform 1 0 8928 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_102
timestamp 1677580104
transform 1 0 10368 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_104
timestamp 1677579658
transform 1 0 10560 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_114
timestamp 1677580104
transform 1 0 11520 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_116
timestamp 1677579658
transform 1 0 11712 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_130
timestamp 1679581782
transform 1 0 13056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_137
timestamp 1679581782
transform 1 0 13728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_0
timestamp 1679577901
transform 1 0 576 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_4
timestamp 1677579658
transform 1 0 960 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_32
timestamp 1679577901
transform 1 0 3648 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_72
timestamp 1677580104
transform 1 0 7488 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_74
timestamp 1677579658
transform 1 0 7680 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_88
timestamp 1677579658
transform 1 0 9024 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_120
timestamp 1679581782
transform 1 0 12096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_127
timestamp 1679581782
transform 1 0 12768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_134
timestamp 1679581782
transform 1 0 13440 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_141
timestamp 1677580104
transform 1 0 14112 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_143
timestamp 1677579658
transform 1 0 14304 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 576 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_7
timestamp 1677580104
transform 1 0 1248 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_9
timestamp 1677579658
transform 1 0 1440 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_14
timestamp 1677580104
transform 1 0 1920 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_86
timestamp 1677579658
transform 1 0 8832 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_95
timestamp 1679577901
transform 1 0 9696 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_4  FILLER_9_103
timestamp 1679577901
transform 1 0 10464 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_107
timestamp 1677579658
transform 1 0 10848 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_116
timestamp 1677579658
transform 1 0 11712 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 1248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 1920 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_21
timestamp 1677580104
transform 1 0 2592 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_23
timestamp 1677579658
transform 1 0 2784 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_81
timestamp 1679577901
transform 1 0 8352 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_85
timestamp 1677580104
transform 1 0 8736 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_10_94
timestamp 1679577901
transform 1 0 9600 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_98
timestamp 1677580104
transform 1 0 9984 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_105
timestamp 1677580104
transform 1 0 10656 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1679581782
transform 1 0 1248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1679581782
transform 1 0 1920 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_21
timestamp 1677580104
transform 1 0 2592 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_23
timestamp 1677579658
transform 1 0 2784 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_36
timestamp 1679581782
transform 1 0 4032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_43
timestamp 1679577901
transform 1 0 4704 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_47
timestamp 1677579658
transform 1 0 5088 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_80
timestamp 1677580104
transform 1 0 8256 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_109
timestamp 1677579658
transform 1 0 11040 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_143
timestamp 1677579658
transform 1 0 14304 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_0
timestamp 1679581782
transform 1 0 576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_7
timestamp 1679581782
transform 1 0 1248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_14
timestamp 1679581782
transform 1 0 1920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_21
timestamp 1679581782
transform 1 0 2592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_28
timestamp 1679581782
transform 1 0 3264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_35
timestamp 1679577901
transform 1 0 3936 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_39
timestamp 1677579658
transform 1 0 4320 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_57
timestamp 1677580104
transform 1 0 6048 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_63
timestamp 1677580104
transform 1 0 6624 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_73
timestamp 1679581782
transform 1 0 7584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_80
timestamp 1679581782
transform 1 0 8256 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_92
timestamp 1677579658
transform 1 0 9408 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_103
timestamp 1677580104
transform 1 0 10464 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_12_135
timestamp 1679581782
transform 1 0 13536 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_142
timestamp 1677580104
transform 1 0 14208 0 1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_4
timestamp 1679581782
transform 1 0 960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_11
timestamp 1679577901
transform 1 0 1632 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_15
timestamp 1677579658
transform 1 0 2016 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_70
timestamp 1677579658
transform 1 0 7296 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_124
timestamp 1679581782
transform 1 0 12480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_131
timestamp 1679581782
transform 1 0 13152 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_138
timestamp 1677580104
transform 1 0 13824 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_27
timestamp 1677579658
transform 1 0 3168 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_55
timestamp 1679577901
transform 1 0 5856 0 1 11340
box -48 -56 432 834
use sg13g2_decap_4  FILLER_15_0
timestamp 1679577901
transform 1 0 576 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_4
timestamp 1677579658
transform 1 0 960 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_9
timestamp 1679581782
transform 1 0 1440 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_16
timestamp 1677580104
transform 1 0 2112 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_31
timestamp 1677579658
transform 1 0 3552 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_59
timestamp 1679577901
transform 1 0 6240 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_63
timestamp 1677579658
transform 1 0 6624 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_68
timestamp 1677579658
transform 1 0 7104 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_99
timestamp 1677580104
transform 1 0 10080 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_132
timestamp 1679581782
transform 1 0 13248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_15_139
timestamp 1679577901
transform 1 0 13920 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_143
timestamp 1677579658
transform 1 0 14304 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_0
timestamp 1679581782
transform 1 0 576 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_7
timestamp 1679581782
transform 1 0 1248 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_14
timestamp 1679581782
transform 1 0 1920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_21
timestamp 1679581782
transform 1 0 2592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_28
timestamp 1679581782
transform 1 0 3264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_35
timestamp 1679581782
transform 1 0 3936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_42
timestamp 1679577901
transform 1 0 4608 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_46
timestamp 1677580104
transform 1 0 4992 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_52
timestamp 1679581782
transform 1 0 5568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_59
timestamp 1679577901
transform 1 0 6240 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_81
timestamp 1677580104
transform 1 0 8352 0 1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_90
timestamp 1677580104
transform 1 0 9216 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_114
timestamp 1677579658
transform 1 0 11520 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_124
timestamp 1679581782
transform 1 0 12480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_131
timestamp 1679581782
transform 1 0 13152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_138
timestamp 1679577901
transform 1 0 13824 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_142
timestamp 1677580104
transform 1 0 14208 0 1 12852
box -48 -56 240 834
use sg13g2_dlygate4sd3_1  hold1
timestamp 1677672058
transform -1 0 3552 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold2
timestamp 1677672058
transform -1 0 4896 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold3
timestamp 1677672058
transform -1 0 6240 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold4
timestamp 1677672058
transform 1 0 9984 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold5
timestamp 1677672058
transform -1 0 3456 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold6
timestamp 1677672058
transform -1 0 10176 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold7
timestamp 1677672058
transform -1 0 8640 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold8
timestamp 1677672058
transform -1 0 6048 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold9
timestamp 1677672058
transform -1 0 4896 0 1 756
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold10
timestamp 1677672058
transform -1 0 7584 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1677672058
transform -1 0 6624 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1677672058
transform -1 0 9312 0 1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1677672058
transform -1 0 7776 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1677672058
transform -1 0 7488 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1677672058
transform -1 0 13536 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1677672058
transform 1 0 10848 0 1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1677672058
transform -1 0 13056 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677672058
transform -1 0 12192 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677672058
transform -1 0 11328 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677672058
transform 1 0 4992 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677672058
transform -1 0 6720 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677672058
transform -1 0 4320 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677672058
transform -1 0 2976 0 -1 8316
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677672058
transform 1 0 6048 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677672058
transform 1 0 7488 0 1 2268
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677672058
transform -1 0 5760 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677672058
transform -1 0 4896 0 1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677672058
transform -1 0 13920 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677672058
transform -1 0 12672 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1677672058
transform -1 0 10176 0 1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1677672058
transform 1 0 8352 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold32
timestamp 1677672058
transform -1 0 9216 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold33
timestamp 1677672058
transform -1 0 8352 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold34
timestamp 1677672058
transform -1 0 11520 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold35
timestamp 1677672058
transform -1 0 9984 0 -1 6804
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold36
timestamp 1677672058
transform -1 0 12480 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold37
timestamp 1677672058
transform -1 0 11712 0 -1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold38
timestamp 1677672058
transform -1 0 10272 0 1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold39
timestamp 1677672058
transform -1 0 10080 0 -1 12852
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold40
timestamp 1677672058
transform -1 0 9792 0 1 11340
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold41
timestamp 1677672058
transform -1 0 5280 0 -1 5292
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold42
timestamp 1677672058
transform -1 0 13440 0 -1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold43
timestamp 1677672058
transform -1 0 11520 0 1 9828
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold44
timestamp 1677672058
transform -1 0 10176 0 -1 3780
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold45
timestamp 1677672058
transform -1 0 6240 0 1 3780
box -48 -56 912 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output2
timestamp 1676381911
transform 1 0 14016 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output3
timestamp 1676381911
transform 1 0 14016 0 -1 11340
box -48 -56 432 834
<< labels >>
flabel metal4 s 4316 712 4756 13652 0 FreeSans 2560 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 532 4496 14444 4936 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3076 712 3516 13652 0 FreeSans 2560 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 532 3256 14444 3696 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 14920 3740 15000 3820 0 FreeSans 320 0 0 0 env_bit
port 3 nsew signal output
flabel metal3 s 14920 11132 15000 11212 0 FreeSans 320 0 0 0 env_valid
port 4 nsew signal output
flabel metal3 s 0 11132 80 11212 0 FreeSans 320 0 0 0 spad_hit_async
port 5 nsew signal input
rlabel metal1 7488 12852 7488 12852 0 VGND
rlabel metal1 7488 13608 7488 13608 0 VPWR
rlabel metal2 4800 11676 4800 11676 0 _000_
rlabel metal2 5664 9408 5664 9408 0 _001_
rlabel metal2 11136 8400 11136 8400 0 _002_
rlabel metal3 6816 11676 6816 11676 0 _003_
rlabel metal2 9312 11004 9312 11004 0 _004_
rlabel metal2 10464 9660 10464 9660 0 _005_
rlabel metal3 8976 8820 8976 8820 0 _006_
rlabel metal3 1296 4368 1296 4368 0 _007_
rlabel metal2 2016 3822 2016 3822 0 _008_
rlabel metal3 4494 3528 4494 3528 0 _009_
rlabel metal2 4800 1134 4800 1134 0 _010_
rlabel metal3 7104 2604 7104 2604 0 _011_
rlabel metal2 8448 3486 8448 3486 0 _012_
rlabel metal2 8496 2604 8496 2604 0 _013_
rlabel metal3 8064 7140 8064 7140 0 _014_
rlabel metal3 11712 3612 11712 3612 0 _015_
rlabel metal3 10800 4116 10800 4116 0 _016_
rlabel metal2 9888 6720 9888 6720 0 _017_
rlabel metal2 5184 6132 5184 6132 0 _018_
rlabel metal3 5136 7140 5136 7140 0 _019_
rlabel metal2 3024 8148 3024 8148 0 _020_
rlabel metal2 2880 8694 2880 8694 0 _021_
rlabel metal2 5952 6888 5952 6888 0 _022_
rlabel metal3 13392 8064 13392 8064 0 _023_
rlabel metal3 3840 7980 3840 7980 0 _024_
rlabel metal3 7632 4956 7632 4956 0 _025_
rlabel metal2 5472 8904 5472 8904 0 _026_
rlabel metal2 4800 3276 4800 3276 0 _027_
rlabel metal2 6432 3360 6432 3360 0 _028_
rlabel metal2 7008 3809 7008 3809 0 _029_
rlabel metal2 6720 4998 6720 4998 0 _030_
rlabel metal3 9744 3444 9744 3444 0 _031_
rlabel metal2 6816 4914 6816 4914 0 _032_
rlabel metal3 7344 5628 7344 5628 0 _033_
rlabel metal3 8160 7056 8160 7056 0 _034_
rlabel metal2 5664 5670 5664 5670 0 _035_
rlabel metal2 4512 6090 4512 6090 0 _036_
rlabel metal2 6144 5880 6144 5880 0 _037_
rlabel metal2 12048 10164 12048 10164 0 _038_
rlabel metal2 11760 10164 11760 10164 0 _039_
rlabel metal2 11424 9450 11424 9450 0 _040_
rlabel metal2 13536 9534 13536 9534 0 _041_
rlabel metal3 12432 7980 12432 7980 0 _042_
rlabel metal2 7680 12936 7680 12936 0 _043_
rlabel metal2 9984 12558 9984 12558 0 _044_
rlabel metal2 9072 13104 9072 13104 0 _045_
rlabel metal2 11568 11004 11568 11004 0 _046_
rlabel metal2 10272 10206 10272 10206 0 _047_
rlabel metal2 10176 10122 10176 10122 0 _048_
rlabel metal2 9504 9324 9504 9324 0 _049_
rlabel metal2 6144 4872 6144 4872 0 _050_
rlabel metal2 7968 4032 7968 4032 0 _051_
rlabel metal2 10848 3822 10848 3822 0 _052_
rlabel metal2 7680 5208 7680 5208 0 _053_
rlabel metal3 1182 3780 1182 3780 0 clk
rlabel metal2 4944 8064 4944 8064 0 clknet_0_clk
rlabel metal2 3264 2562 3264 2562 0 clknet_2_0__leaf_clk
rlabel metal3 2688 11004 2688 11004 0 clknet_2_1__leaf_clk
rlabel metal3 9984 4788 9984 4788 0 clknet_2_2__leaf_clk
rlabel metal2 13056 8316 13056 8316 0 clknet_2_3__leaf_clk
rlabel metal3 14630 3780 14630 3780 0 env_bit
rlabel metal3 14630 11172 14630 11172 0 env_valid
rlabel metal2 672 11382 672 11382 0 net1
rlabel metal2 2496 3864 2496 3864 0 net10
rlabel metal2 2112 3444 2112 3444 0 net11
rlabel metal2 1344 5376 1344 5376 0 net12
rlabel metal2 13968 9324 13968 9324 0 net13
rlabel metal2 9024 9156 9024 9156 0 net14
rlabel metal3 12624 12348 12624 12348 0 net15
rlabel metal2 11232 12936 11232 12936 0 net16
rlabel metal2 6240 8736 6240 8736 0 net17
rlabel metal2 6912 12180 6912 12180 0 net18
rlabel metal2 1584 7812 1584 7812 0 net19
rlabel metal2 14160 8652 14160 8652 0 net2
rlabel metal2 6768 11676 6768 11676 0 net20
rlabel metal2 3744 8988 3744 8988 0 net21
rlabel metal2 3072 5796 3072 5796 0 net22
rlabel metal2 6864 10332 6864 10332 0 net23
rlabel metal2 10080 6720 10080 6720 0 net24
rlabel metal3 11376 7308 11376 7308 0 net25
rlabel metal2 12528 4956 12528 4956 0 net26
rlabel metal2 8304 4284 8304 4284 0 net27
rlabel metal3 9552 3276 9552 3276 0 net28
rlabel metal2 9408 1596 9408 1596 0 net29
rlabel metal2 14112 11214 14112 11214 0 net3
rlabel metal3 7536 1260 7536 1260 0 net30
rlabel metal2 5232 13356 5232 13356 0 net31
rlabel metal2 2208 11676 2208 11676 0 net32
rlabel metal2 4128 11970 4128 11970 0 net33
rlabel metal2 5376 12516 5376 12516 0 net34
rlabel metal2 8976 10164 8976 10164 0 net35
rlabel metal3 2208 4116 2208 4116 0 net36
rlabel metal3 8352 5880 8352 5880 0 net37
rlabel metal2 7872 6006 7872 6006 0 net38
rlabel metal2 5280 2898 5280 2898 0 net39
rlabel metal2 3648 3108 3648 3108 0 net4
rlabel metal3 3552 1260 3552 1260 0 net40
rlabel metal2 5616 8652 5616 8652 0 net41
rlabel metal2 5856 7980 5856 7980 0 net42
rlabel metal2 8592 5880 8592 5880 0 net43
rlabel metal2 5184 5376 5184 5376 0 net44
rlabel metal2 6432 6594 6432 6594 0 net45
rlabel metal2 12192 9786 12192 9786 0 net46
rlabel metal2 11712 8652 11712 8652 0 net47
rlabel metal3 12096 3444 12096 3444 0 net48
rlabel metal2 11424 4746 11424 4746 0 net49
rlabel metal2 6144 9912 6144 9912 0 net5
rlabel metal2 10560 4956 10560 4956 0 net50
rlabel metal3 5376 5460 5376 5460 0 net51
rlabel metal2 5952 8904 5952 8904 0 net52
rlabel metal2 3552 8820 3552 8820 0 net53
rlabel metal2 1152 7434 1152 7434 0 net54
rlabel metal2 6240 2982 6240 2982 0 net55
rlabel metal2 8304 2016 8304 2016 0 net56
rlabel metal3 5328 5628 5328 5628 0 net57
rlabel metal3 3408 6468 3408 6468 0 net58
rlabel metal2 12096 3696 12096 3696 0 net59
rlabel metal2 12240 8652 12240 8652 0 net6
rlabel metal2 11904 5628 11904 5628 0 net60
rlabel metal2 7680 3486 7680 3486 0 net61
rlabel metal2 8592 2016 8592 2016 0 net62
rlabel metal2 7872 12684 7872 12684 0 net63
rlabel metal3 7440 12516 7440 12516 0 net64
rlabel metal3 9840 7140 9840 7140 0 net65
rlabel metal2 9216 6846 9216 6846 0 net66
rlabel metal3 11376 13020 11376 13020 0 net67
rlabel metal2 10368 9030 10368 9030 0 net68
rlabel metal3 8112 13188 8112 13188 0 net69
rlabel metal2 1104 12348 1104 12348 0 net7
rlabel metal2 9216 11214 9216 11214 0 net70
rlabel metal3 8256 11088 8256 11088 0 net71
rlabel metal3 4752 4704 4752 4704 0 net72
rlabel metal3 12384 9492 12384 9492 0 net73
rlabel metal3 10560 10164 10560 10164 0 net74
rlabel metal2 7200 3402 7200 3402 0 net75
rlabel metal2 5376 4032 5376 4032 0 net76
rlabel metal2 2592 11676 2592 11676 0 net8
rlabel metal2 3744 12012 3744 12012 0 net9
rlabel metal3 11712 9492 11712 9492 0 prev2_bit
rlabel metal3 9408 11844 9408 11844 0 pulse_cnt\[0\]
rlabel metal2 10176 12432 10176 12432 0 pulse_cnt\[1\]
rlabel metal3 12432 12264 12432 12264 0 pulse_cnt\[2\]
rlabel metal3 11232 10164 11232 10164 0 pulse_cnt\[3\]
rlabel metal2 7200 12180 7200 12180 0 rise_spad
rlabel metal2 3024 11928 3024 11928 0 s0
rlabel metal2 4752 10920 4752 10920 0 s1
rlabel metal2 5760 12222 5760 12222 0 s1_d
rlabel metal3 462 11172 462 11172 0 spad_hit_async
rlabel metal2 3456 4116 3456 4116 0 win_cnt\[0\]
rlabel metal3 9792 5964 9792 5964 0 win_cnt\[10\]
rlabel metal3 9024 5628 9024 5628 0 win_cnt\[11\]
rlabel metal3 5424 6216 5424 6216 0 win_cnt\[12\]
rlabel metal2 5088 8232 5088 8232 0 win_cnt\[13\]
rlabel metal2 3552 6846 3552 6846 0 win_cnt\[14\]
rlabel metal3 7872 7980 7872 7980 0 win_cnt\[15\]
rlabel metal2 5472 3381 5472 3381 0 win_cnt\[1\]
rlabel metal2 5664 3780 5664 3780 0 win_cnt\[2\]
rlabel metal2 5568 2352 5568 2352 0 win_cnt\[3\]
rlabel metal2 6000 2100 6000 2100 0 win_cnt\[4\]
rlabel metal3 10464 2100 10464 2100 0 win_cnt\[5\]
rlabel metal3 10464 2856 10464 2856 0 win_cnt\[6\]
rlabel metal2 10272 5250 10272 5250 0 win_cnt\[7\]
rlabel metal2 13824 3948 13824 3948 0 win_cnt\[8\]
rlabel metal2 12960 4788 12960 4788 0 win_cnt\[9\]
rlabel metal2 8160 9786 8160 9786 0 win_rollover
<< properties >>
string FIXED_BBOX 0 0 15000 15000
<< end >>
